magic
tech scmos
timestamp 951727448
<< pwell >>
rect 0 0 40 32
<< nwell >>
rect 0 32 40 64
<< polysilicon >>
rect 11 56 29 58
rect 11 52 13 56
rect 15 52 17 54
rect 23 52 25 54
rect 27 52 29 56
rect 11 24 13 44
rect 15 43 17 44
rect 23 43 25 44
rect 15 41 25 43
rect 27 42 29 44
rect 23 37 25 41
rect 19 24 21 37
rect 11 10 13 12
rect 19 10 21 12
<< ndiffusion >>
rect 10 12 11 24
rect 13 12 14 24
rect 18 12 19 24
rect 21 12 22 24
<< pdiffusion >>
rect 10 44 11 52
rect 13 44 15 52
rect 17 44 18 52
rect 22 44 23 52
rect 25 44 27 52
rect 29 44 30 52
<< metal1 >>
rect 0 56 6 60
rect 10 56 30 60
rect 34 56 40 60
rect 6 52 10 56
rect 30 52 34 56
rect 7 32 10 33
rect 14 30 18 47
rect 22 32 25 33
rect 14 24 18 26
rect 6 8 10 12
rect 22 8 26 12
rect 0 4 6 8
rect 10 4 22 8
rect 26 4 30 8
rect 34 4 40 8
<< ntransistor >>
rect 11 12 13 24
rect 19 12 21 24
<< ptransistor >>
rect 11 44 13 52
rect 15 44 17 52
rect 23 44 25 52
rect 27 44 29 52
<< polycontact >>
rect 7 33 11 37
rect 21 33 25 37
<< ndcontact >>
rect 6 12 10 24
rect 14 12 18 24
rect 22 12 26 24
<< pdcontact >>
rect 6 44 10 52
rect 18 44 22 52
rect 30 44 34 52
<< m2contact >>
rect 6 28 10 32
rect 14 26 18 30
rect 22 28 26 32
<< psubstratepcontact >>
rect 6 4 10 8
rect 22 4 26 8
rect 30 4 34 8
<< nsubstratencontact >>
rect 6 56 10 60
rect 30 56 34 60
<< labels >>
rlabel metal1 4 6 4 6 6 GND
rlabel metal1 36 6 36 6 6 GND
rlabel metal1 4 58 4 58 6 Vdd
rlabel metal1 36 58 36 58 6 Vdd
rlabel m2contact 8 30 8 30 6 In1
rlabel m2contact 16 28 16 28 6 Out_b
rlabel m2contact 24 30 24 30 6 In0
<< end >>
