magic
tech scmos
timestamp 951209823
<< nwell >>
rect 122 -26 209 37
<< polysilicon >>
rect 53 25 64 27
rect 69 25 71 27
rect 53 20 55 25
rect 90 20 124 22
rect 73 15 75 17
rect 83 15 89 17
rect 128 14 131 16
rect 147 14 149 16
rect 156 15 158 17
rect 168 15 173 17
rect 48 7 50 9
rect 55 8 58 9
rect 185 8 188 9
rect 55 7 72 8
rect 56 6 68 7
rect 164 7 188 8
rect 198 7 200 9
rect 48 -1 50 1
rect 55 0 58 1
rect 168 6 187 7
rect 185 0 188 1
rect 55 -1 59 0
rect 56 -2 59 -1
rect 64 -2 77 0
rect 93 -2 124 0
rect 156 -2 174 0
rect 184 -1 188 0
rect 198 -1 200 1
rect 184 -2 187 -1
rect 48 -10 50 -8
rect 55 -10 59 -8
rect 64 -10 68 -8
rect 73 -10 77 -8
rect 93 -10 96 -8
rect 100 -10 124 -8
rect 156 -10 160 -8
rect 170 -10 174 -8
rect 184 -10 188 -8
rect 198 -10 200 -8
rect 48 -18 50 -16
rect 55 -18 59 -16
rect 64 -18 68 -16
rect 73 -18 77 -16
rect 93 -18 117 -16
rect 121 -18 124 -16
rect 156 -18 160 -16
rect 170 -18 174 -16
rect 184 -18 188 -16
rect 198 -18 200 -16
<< ndiffusion >>
rect 64 27 69 28
rect 64 24 69 25
rect 75 17 83 18
rect 75 14 83 15
rect 50 9 55 10
rect 50 6 55 7
rect 50 1 55 2
rect 59 0 64 1
rect 77 0 93 1
rect 50 -2 55 -1
rect 44 -7 55 -2
rect 50 -8 55 -7
rect 59 -8 64 -2
rect 77 -3 93 -2
rect 68 -8 73 -7
rect 77 -8 93 -7
rect 50 -11 55 -10
rect 50 -16 55 -15
rect 59 -16 64 -10
rect 68 -16 73 -10
rect 77 -11 93 -10
rect 86 -15 93 -11
rect 77 -16 93 -15
rect 50 -19 55 -18
rect 59 -19 64 -18
rect 68 -19 73 -18
rect 77 -19 93 -18
<< pdiffusion >>
rect 158 17 168 18
rect 131 16 147 17
rect 158 14 168 15
rect 131 13 147 14
rect 188 9 198 10
rect 188 6 198 7
rect 124 0 156 1
rect 188 1 198 2
rect 174 0 184 1
rect 188 -2 198 -1
rect 124 -3 156 -2
rect 124 -8 156 -7
rect 160 -8 170 -7
rect 174 -8 184 -2
rect 188 -7 201 -2
rect 188 -8 198 -7
rect 124 -11 156 -10
rect 124 -15 131 -11
rect 124 -16 156 -15
rect 160 -16 170 -10
rect 174 -16 184 -10
rect 188 -11 198 -10
rect 188 -16 198 -15
rect 124 -19 156 -18
rect 160 -19 170 -18
rect 174 -19 184 -18
rect 188 -19 198 -18
<< metal1 >>
rect 69 28 97 32
rect 93 27 97 28
rect 44 24 61 26
rect 44 23 64 24
rect 44 -7 47 23
rect 58 20 64 23
rect 69 20 70 24
rect 55 16 56 17
rect 51 14 56 16
rect 55 13 56 14
rect 60 13 63 17
rect 40 -11 44 -7
rect 51 -11 55 2
rect 59 5 63 13
rect 67 13 70 20
rect 83 18 86 24
rect 67 10 75 13
rect 89 10 93 13
rect 89 5 93 6
rect 72 3 77 5
rect 68 1 77 3
rect 68 -3 72 1
rect 68 -15 77 -11
rect 40 -19 44 -15
rect 68 -19 72 -15
rect 89 -19 93 -7
rect 96 -11 100 -10
rect 103 -18 106 37
rect 40 -23 50 -19
rect 55 -23 59 -19
rect 64 -23 68 -19
rect 111 -27 114 24
rect 128 21 147 23
rect 128 20 131 21
rect 150 14 153 33
rect 158 22 169 26
rect 124 10 128 13
rect 150 12 158 14
rect 147 10 158 12
rect 177 13 178 17
rect 182 14 194 17
rect 147 9 153 10
rect 124 5 128 6
rect 156 3 164 5
rect 176 5 182 13
rect 156 1 168 3
rect 162 -3 168 1
rect 117 -16 121 -15
rect 124 -19 128 -7
rect 190 -11 196 2
rect 201 -2 205 33
rect 156 -15 168 -11
rect 162 -19 168 -15
rect 201 -19 205 -7
rect 170 -23 174 -19
rect 184 -23 188 -19
rect 198 -23 202 -19
rect 207 -23 209 -19
<< metal2 >>
rect 40 33 150 37
rect 154 33 201 37
rect 205 33 209 37
rect 40 32 209 33
rect 40 31 208 32
rect 40 23 93 26
rect 97 23 169 26
rect 40 22 169 23
rect 173 22 209 26
rect 56 17 182 18
rect 60 14 178 17
rect 93 6 124 10
rect 40 0 55 1
rect 40 -4 209 0
rect 40 -14 96 -11
rect 121 -14 209 -11
rect 40 -23 209 -21
rect 44 -27 209 -23
<< ntransistor >>
rect 64 25 69 27
rect 75 15 83 17
rect 50 7 55 9
rect 50 -1 55 1
rect 59 -2 64 0
rect 77 -2 93 0
rect 50 -10 55 -8
rect 59 -10 64 -8
rect 68 -10 73 -8
rect 77 -10 93 -8
rect 50 -18 55 -16
rect 59 -18 64 -16
rect 68 -18 73 -16
rect 77 -18 93 -16
<< ptransistor >>
rect 131 14 147 16
rect 158 15 168 17
rect 188 7 198 9
rect 124 -2 156 0
rect 174 -2 184 0
rect 188 -1 198 1
rect 124 -10 156 -8
rect 160 -10 170 -8
rect 174 -10 184 -8
rect 188 -10 198 -8
rect 124 -18 156 -16
rect 160 -18 170 -16
rect 174 -18 184 -16
rect 188 -18 198 -16
<< polycontact >>
rect 51 16 55 20
rect 86 20 90 24
rect 124 20 128 24
rect 89 13 93 17
rect 124 13 128 17
rect 173 13 177 17
rect 68 3 72 7
rect 164 3 168 7
rect 96 -10 100 -6
rect 117 -20 121 -16
<< ndcontact >>
rect 64 28 69 32
rect 64 20 69 24
rect 75 18 83 22
rect 50 10 55 14
rect 75 10 83 14
rect 50 2 55 6
rect 59 1 64 5
rect 77 1 93 5
rect 40 -7 44 -2
rect 68 -7 73 -3
rect 77 -7 93 -3
rect 50 -15 55 -11
rect 77 -15 86 -11
rect 50 -23 55 -19
rect 59 -23 64 -19
rect 68 -23 73 -19
rect 77 -23 93 -19
<< pdcontact >>
rect 131 17 147 21
rect 158 18 168 22
rect 131 9 147 13
rect 158 10 168 14
rect 188 10 198 14
rect 124 1 156 5
rect 174 1 184 5
rect 188 2 198 6
rect 124 -7 156 -3
rect 160 -7 170 -3
rect 201 -7 205 -2
rect 131 -15 156 -11
rect 188 -15 198 -11
rect 124 -23 156 -19
rect 160 -23 170 -19
rect 174 -23 184 -19
rect 188 -23 198 -19
<< m2contact >>
rect 56 13 60 17
rect 93 23 97 27
rect 89 6 93 10
rect 96 -15 100 -11
rect 150 33 154 37
rect 201 33 205 37
rect 40 -27 44 -23
rect 169 22 173 26
rect 124 6 128 10
rect 178 13 182 17
rect 117 -15 121 -11
<< psubstratepcontact >>
rect 40 -15 44 -11
<< nsubstratencontact >>
rect 202 -23 207 -19
<< labels >>
rlabel polysilicon 99 20 99 20 1 Cout
rlabel polysilicon 98 -1 98 -1 1 Cin
rlabel metal2 47 -25 47 -25 1 Gnd
rlabel metal2 47 -13 47 -13 1 A
rlabel metal2 47 34 47 34 5 Vdd
rlabel metal2 167 16 167 16 1 Sum_b
rlabel metal2 207 -13 207 -13 7 B
rlabel metal2 207 -2 207 -2 7 Random
rlabel metal2 207 24 207 24 7 Sum
<< end >>
