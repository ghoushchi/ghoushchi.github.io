magic
tech scmos
timestamp 950486748
<< metal1 >>
rect 67 168 219 320
rect 19 115 237 117
rect 19 111 25 115
rect 29 111 30 115
rect 34 111 35 115
rect 39 113 237 115
rect 241 113 242 117
rect 246 113 247 117
rect 251 113 261 117
rect 39 112 261 113
rect 39 111 237 112
rect 19 110 237 111
rect 19 106 25 110
rect 29 106 30 110
rect 34 106 35 110
rect 39 108 237 110
rect 241 108 242 112
rect 246 108 247 112
rect 251 108 261 112
rect 39 106 261 108
rect 19 105 261 106
rect 11 101 12 105
rect 260 101 261 105
rect 19 99 261 101
rect 19 96 237 99
rect 19 92 25 96
rect 29 92 30 96
rect 34 92 35 96
rect 39 95 237 96
rect 241 95 242 99
rect 246 95 247 99
rect 251 95 261 99
rect 39 94 261 95
rect 39 92 237 94
rect 19 91 237 92
rect 19 87 25 91
rect 29 87 30 91
rect 34 87 35 91
rect 39 90 237 91
rect 241 90 242 94
rect 246 90 247 94
rect 251 90 261 94
rect 39 89 261 90
rect 39 87 237 89
rect 19 86 237 87
rect 19 82 25 86
rect 29 82 30 86
rect 34 82 35 86
rect 39 85 237 86
rect 241 85 242 89
rect 246 85 247 89
rect 251 85 261 89
rect 39 84 261 85
rect 39 82 237 84
rect 19 81 237 82
rect 19 77 25 81
rect 29 77 30 81
rect 34 77 35 81
rect 39 80 237 81
rect 241 80 242 84
rect 246 80 247 84
rect 251 80 261 84
rect 39 79 261 80
rect 39 77 237 79
rect 19 76 237 77
rect 19 72 25 76
rect 29 72 30 76
rect 34 72 35 76
rect 39 75 237 76
rect 241 75 242 79
rect 246 75 247 79
rect 251 75 261 79
rect 39 74 261 75
rect 39 72 237 74
rect 19 70 237 72
rect 241 70 242 74
rect 246 70 247 74
rect 251 70 261 74
rect 28 37 29 41
rect 33 37 34 41
rect 24 36 38 37
rect 28 32 29 36
rect 33 32 34 36
rect 24 31 38 32
rect 28 27 29 31
rect 33 27 34 31
rect 25 17 37 27
rect 52 5 236 6
rect 68 1 72 5
rect 76 1 80 5
rect 84 1 88 5
rect 92 1 96 5
rect 100 1 104 5
rect 108 1 112 5
rect 116 1 120 5
rect 124 1 128 5
rect 132 1 136 5
rect 140 1 144 5
rect 148 1 152 5
rect 156 1 160 5
rect 164 1 168 5
rect 172 1 176 5
rect 180 1 184 5
rect 188 1 192 5
rect 196 1 200 5
rect 204 1 208 5
rect 212 1 216 5
rect 220 1 224 5
rect 52 0 236 1
<< metal2 >>
rect 68 315 218 319
rect 68 173 72 315
rect 214 173 218 315
rect 68 169 218 173
rect 0 115 39 116
rect 0 111 25 115
rect 29 111 30 115
rect 34 111 35 115
rect 0 110 39 111
rect 0 106 25 110
rect 29 106 30 110
rect 34 106 35 110
rect 0 96 39 106
rect 0 92 25 96
rect 29 92 30 96
rect 34 92 35 96
rect 0 91 39 92
rect 0 87 25 91
rect 29 87 30 91
rect 34 87 35 91
rect 0 86 39 87
rect 0 82 25 86
rect 29 82 30 86
rect 34 82 35 86
rect 0 81 39 82
rect 0 77 25 81
rect 29 77 30 81
rect 34 77 35 81
rect 0 76 39 77
rect 0 72 25 76
rect 29 72 30 76
rect 34 72 35 76
rect 0 70 39 72
rect 68 58 219 169
rect 241 113 242 117
rect 246 113 247 117
rect 251 113 285 116
rect 237 112 285 113
rect 241 108 242 112
rect 246 108 247 112
rect 251 108 285 112
rect 237 99 285 108
rect 241 95 242 99
rect 246 95 247 99
rect 251 95 285 99
rect 237 94 285 95
rect 241 90 242 94
rect 246 90 247 94
rect 251 90 285 94
rect 237 89 285 90
rect 241 85 242 89
rect 246 85 247 89
rect 251 85 285 89
rect 237 84 285 85
rect 241 80 242 84
rect 246 80 247 84
rect 251 80 285 84
rect 237 79 285 80
rect 241 75 242 79
rect 246 75 247 79
rect 251 75 285 79
rect 237 74 285 75
rect 241 70 242 74
rect 246 70 247 74
rect 251 70 285 74
rect 0 41 285 58
rect 0 37 24 41
rect 28 37 29 41
rect 33 37 34 41
rect 38 37 285 41
rect 0 36 285 37
rect 0 32 24 36
rect 28 32 29 36
rect 33 32 34 36
rect 38 32 285 36
rect 0 31 285 32
rect 0 27 24 31
rect 28 27 29 31
rect 33 27 34 31
rect 38 27 285 31
rect 0 10 285 27
rect 0 5 60 6
rect 0 1 40 5
rect 44 1 48 5
rect 52 1 56 5
rect 0 0 60 1
rect 68 0 219 10
rect 227 5 285 6
rect 227 1 228 5
rect 232 1 236 5
rect 240 1 244 5
rect 248 1 252 5
rect 256 1 260 5
rect 264 1 268 5
rect 272 1 285 5
rect 227 0 285 1
<< m2contact >>
rect 25 111 29 115
rect 30 111 34 115
rect 35 111 39 115
rect 237 113 241 117
rect 242 113 246 117
rect 247 113 251 117
rect 25 106 29 110
rect 30 106 34 110
rect 35 106 39 110
rect 237 108 241 112
rect 242 108 246 112
rect 247 108 251 112
rect 25 92 29 96
rect 30 92 34 96
rect 35 92 39 96
rect 237 95 241 99
rect 242 95 246 99
rect 247 95 251 99
rect 25 87 29 91
rect 30 87 34 91
rect 35 87 39 91
rect 237 90 241 94
rect 242 90 246 94
rect 247 90 251 94
rect 25 82 29 86
rect 30 82 34 86
rect 35 82 39 86
rect 237 85 241 89
rect 242 85 246 89
rect 247 85 251 89
rect 25 77 29 81
rect 30 77 34 81
rect 35 77 39 81
rect 237 80 241 84
rect 242 80 246 84
rect 247 80 251 84
rect 25 72 29 76
rect 30 72 34 76
rect 35 72 39 76
rect 237 75 241 79
rect 242 75 246 79
rect 247 75 251 79
rect 237 70 241 74
rect 242 70 246 74
rect 247 70 251 74
rect 24 37 28 41
rect 29 37 33 41
rect 34 37 38 41
rect 24 32 28 36
rect 29 32 33 36
rect 34 32 38 36
rect 24 27 28 31
rect 29 27 33 31
rect 34 27 38 31
rect 40 1 44 5
rect 48 1 52 5
rect 56 1 60 5
rect 228 1 232 5
rect 236 1 240 5
rect 244 1 248 5
rect 252 1 256 5
rect 260 1 264 5
rect 268 1 272 5
<< psubstratepcontact >>
rect 12 101 260 105
rect 44 1 48 5
rect 52 1 56 5
rect 60 1 68 5
rect 72 1 76 5
rect 80 1 84 5
rect 88 1 92 5
rect 96 1 100 5
rect 104 1 108 5
rect 112 1 116 5
rect 120 1 124 5
rect 128 1 132 5
rect 136 1 140 5
rect 144 1 148 5
rect 152 1 156 5
rect 160 1 164 5
rect 168 1 172 5
rect 176 1 180 5
rect 184 1 188 5
rect 192 1 196 5
rect 200 1 204 5
rect 208 1 212 5
rect 216 1 220 5
rect 224 1 228 5
rect 232 1 236 5
rect 240 1 244 5
rect 248 1 252 5
rect 256 1 260 5
rect 264 1 268 5
rect 272 1 276 5
<< nsubstratencontact >>
rect 18 13 258 17
<< psubstratepdiff >>
rect 4 139 281 141
rect 0 133 285 139
rect 0 105 8 133
rect 131 107 160 133
rect 254 107 285 133
rect 131 105 285 107
rect 0 101 12 105
rect 260 101 285 105
rect 0 100 285 101
rect 43 80 47 100
rect 67 80 74 100
rect 187 80 195 100
rect 43 76 195 80
rect 0 5 285 6
rect 0 1 44 5
rect 48 1 52 5
rect 56 1 60 5
rect 68 1 72 5
rect 76 1 80 5
rect 84 1 88 5
rect 92 1 96 5
rect 100 1 104 5
rect 108 1 112 5
rect 116 1 120 5
rect 124 1 128 5
rect 132 1 136 5
rect 140 1 144 5
rect 148 1 152 5
rect 156 1 160 5
rect 164 1 168 5
rect 172 1 176 5
rect 180 1 184 5
rect 188 1 192 5
rect 196 1 200 5
rect 204 1 208 5
rect 212 1 216 5
rect 220 1 224 5
rect 228 1 232 5
rect 236 1 240 5
rect 244 1 248 5
rect 252 1 256 5
rect 260 1 264 5
rect 268 1 272 5
rect 276 1 285 5
rect 0 0 285 1
<< nsubstratendiff >>
rect 0 52 285 56
rect 0 46 6 52
rect 0 18 7 46
rect 43 18 47 52
rect 67 20 80 52
rect 131 50 141 52
rect 174 51 285 52
rect 174 20 188 51
rect 67 18 188 20
rect 272 18 285 51
rect 0 17 285 18
rect 0 13 18 17
rect 258 13 285 17
rect 0 12 285 13
<< pad >>
rect 72 173 214 315
<< glass >>
rect 78 179 208 309
<< labels >>
rlabel space 0 320 0 320 4 sllu_1988
rlabel space 285 320 285 320 6 mosis_tinychip
rlabel metal1 143 234 143 234 6 pad
rlabel metal2 0 70 0 70 4 {w}tiny12_t
rlabel metal2 0 58 0 58 4 {w}tiny12_b
rlabel metal2 285 70 285 70 6 {e}tiny12_t
rlabel metal2 285 58 285 58 6 {e}tiny12_b
rlabel metal2 143 0 143 0 8 .VDD
rlabel psubstratepdiff 0 100 0 100 4 {w}*
rlabel psubstratepdiff 285 100 285 100 6 {e}*
<< end >>
