magic
tech scmos
timestamp 951985653
<< metal1 >>
rect 1266 722 1269 727
rect 1409 722 1413 726
rect 1445 722 1449 726
rect 1452 722 1456 726
rect 1162 616 1166 707
rect 816 603 819 607
rect 1162 591 1166 612
rect 335 542 338 546
rect 264 481 268 505
rect 444 480 448 507
rect 460 497 464 529
rect 715 497 719 587
rect 452 471 456 492
rect 894 481 898 508
rect 902 497 906 587
rect 1162 555 1166 587
rect 1891 545 1900 659
rect 910 497 914 529
rect 902 473 906 493
rect 952 482 956 487
rect 959 482 963 487
rect 995 482 999 487
rect 1716 433 1720 487
rect 1723 415 1727 487
rect 1730 313 1734 487
rect 1737 295 1741 487
rect 1716 81 1720 219
rect 1723 47 1727 261
rect 1730 25 1734 283
rect 1737 103 1741 197
rect 1744 193 1748 487
rect 1787 482 1791 486
rect 1823 482 1827 486
rect 1830 482 1834 486
rect 1751 175 1755 459
rect 1891 425 1900 539
rect 1924 605 1933 719
rect 1924 484 1933 599
rect 1758 73 1762 381
rect 1765 51 1769 339
rect 1891 305 1900 419
rect 1891 185 1900 299
rect 1891 65 1900 179
rect 1891 -85 1900 59
rect 1903 -12 1907 484
rect 1910 -43 1914 484
rect 1917 -77 1921 484
rect 1924 365 1933 479
rect 1924 245 1933 359
rect 1924 125 1933 239
rect 1924 5 1933 119
<< metal2 >>
rect 1528 719 1924 724
rect 1166 708 1173 711
rect 1336 708 1368 711
rect 1336 688 1360 692
rect 1336 675 1340 688
rect 1364 679 1368 708
rect 1522 677 1531 681
rect 1527 659 1891 665
rect 1336 636 1340 653
rect 1336 632 1360 636
rect 1364 616 1368 646
rect 1522 643 1531 647
rect 1166 613 1173 616
rect 1336 613 1368 616
rect 889 598 1172 604
rect 1527 599 1924 605
rect 719 588 723 591
rect 889 588 902 591
rect 1166 588 1173 591
rect 1336 588 1368 591
rect 1336 568 1360 572
rect 889 551 1162 555
rect 1336 553 1340 568
rect 1364 559 1368 588
rect 1522 557 1531 561
rect 440 539 724 544
rect 886 538 1172 546
rect 1528 539 1891 545
rect 439 529 460 533
rect 890 529 910 533
rect 1336 516 1340 533
rect 1336 512 1360 516
rect 440 493 452 496
rect 464 493 715 497
rect 719 493 723 496
rect 889 493 902 496
rect 1364 496 1368 525
rect 1522 523 1531 527
rect 914 493 1172 496
rect 1338 493 1368 496
rect 440 479 446 484
rect 890 479 896 484
rect 1713 479 1772 484
rect 1857 479 1924 484
rect 441 468 450 471
rect 889 468 900 471
rect 1338 468 1368 471
rect -34 458 -29 462
rect 1 460 20 464
rect 446 463 450 468
rect 896 463 900 468
rect 16 452 20 460
rect 439 459 442 461
rect 438 455 445 459
rect 886 455 895 459
rect 1336 448 1360 452
rect 441 431 447 435
rect 889 431 897 435
rect 1336 434 1340 448
rect 1364 440 1368 468
rect 1755 459 1771 463
rect 1888 460 1935 464
rect 1697 429 1716 433
rect 441 419 445 425
rect 888 419 896 425
rect 1714 419 1772 425
rect 1855 419 1891 425
rect 440 409 447 413
rect 889 409 897 413
rect 1336 396 1340 413
rect 1696 411 1723 415
rect -36 382 -30 386
rect 16 384 20 393
rect 1336 392 1360 396
rect 437 385 444 389
rect 886 385 895 389
rect 1 380 20 384
rect 438 383 441 385
rect 446 376 450 381
rect 896 376 900 381
rect 1364 376 1368 405
rect 1762 381 1773 385
rect 1888 380 1935 384
rect 441 373 450 376
rect 889 373 900 376
rect 1338 373 1368 376
rect 441 359 445 365
rect 889 359 896 365
rect 1714 359 1772 365
rect 1856 359 1924 365
rect 441 348 450 351
rect 890 348 900 351
rect 1338 348 1368 351
rect -34 338 -30 342
rect 1 340 20 344
rect 446 343 450 348
rect 896 343 900 348
rect 16 332 20 340
rect 437 339 441 341
rect 437 335 444 339
rect 886 335 896 339
rect 1336 328 1360 332
rect 441 311 447 315
rect 889 311 897 315
rect 1336 311 1340 328
rect 1364 320 1368 348
rect 1769 339 1773 343
rect 1888 340 1935 344
rect 1696 309 1730 313
rect 441 299 445 305
rect 889 299 897 305
rect 1714 299 1772 305
rect 1855 299 1891 305
rect 441 289 447 293
rect 889 289 897 293
rect 1336 276 1340 293
rect 1696 291 1737 295
rect 1336 272 1360 276
rect -34 262 -30 266
rect 16 264 20 272
rect 1 260 20 264
rect 439 265 444 269
rect 886 265 895 269
rect 439 263 442 265
rect 446 256 450 261
rect 896 256 900 261
rect 1364 256 1368 287
rect 1705 283 1730 287
rect 1727 261 1773 265
rect 1888 260 1935 264
rect 441 253 450 256
rect 889 253 900 256
rect 1335 253 1368 256
rect 441 239 445 245
rect 890 239 896 245
rect 1714 239 1772 245
rect 1856 239 1924 245
rect 441 228 450 231
rect 889 228 900 231
rect 1335 228 1368 231
rect -35 218 -30 222
rect 1 220 20 224
rect 446 223 450 228
rect 896 223 900 228
rect 16 212 20 220
rect 439 218 445 219
rect 437 216 445 218
rect 437 215 444 216
rect 887 215 895 219
rect 1336 208 1360 212
rect 441 191 447 195
rect 890 191 897 195
rect 1336 194 1340 208
rect 1364 200 1368 228
rect 1720 219 1775 223
rect 1888 220 1935 224
rect 1709 197 1737 201
rect 1697 189 1744 193
rect 441 179 445 185
rect 890 179 895 185
rect 1714 179 1772 185
rect 1856 179 1891 185
rect 441 169 447 173
rect 890 169 897 173
rect 1336 156 1340 173
rect 1693 171 1751 175
rect 1336 152 1360 156
rect -34 142 -29 146
rect 16 144 20 152
rect 0 140 20 144
rect 439 145 444 149
rect 887 145 894 149
rect 439 143 442 145
rect 887 143 891 145
rect 446 136 450 141
rect 896 136 900 141
rect 1364 136 1368 167
rect 1709 141 1774 145
rect 1888 140 1935 144
rect 441 133 450 136
rect 889 133 900 136
rect 1335 133 1368 136
rect 441 119 444 125
rect 888 119 895 125
rect 1714 119 1771 125
rect 1856 119 1924 125
rect 441 108 450 111
rect 890 108 900 111
rect 1337 108 1368 111
rect -35 98 -30 102
rect 0 100 20 104
rect 447 103 450 108
rect 896 103 900 108
rect 16 92 20 100
rect 439 99 443 101
rect 439 95 445 99
rect 886 95 895 99
rect 1336 88 1360 92
rect 441 73 447 75
rect 441 71 448 73
rect 890 71 897 75
rect 1336 71 1340 88
rect 1364 77 1368 108
rect 1741 99 1774 103
rect 1888 100 1935 104
rect 1707 77 1716 81
rect 444 69 448 71
rect 1696 69 1758 73
rect 441 59 444 65
rect 890 59 894 65
rect 1714 59 1771 65
rect 1857 59 1891 65
rect 440 49 447 53
rect 890 49 897 53
rect 1696 51 1761 55
rect 1336 36 1340 50
rect 1336 32 1360 36
rect -34 22 -29 26
rect 16 24 20 32
rect 0 20 20 24
rect 438 25 444 29
rect 886 25 895 29
rect 438 23 442 25
rect 448 16 452 17
rect 896 16 900 21
rect 1364 16 1368 47
rect 1710 43 1723 47
rect 1734 21 1775 25
rect 1888 20 1935 24
rect 441 13 452 16
rect 889 13 900 16
rect 1337 13 1368 16
rect 439 0 447 5
rect 890 0 895 5
rect 1713 0 1771 5
rect 1856 0 1924 5
rect -30 -9 1119 -5
rect -30 -17 1067 -13
rect 1115 -14 1119 -9
rect 1384 -16 1903 -12
rect -30 -25 1019 -21
rect 1384 -24 1388 -16
rect 1570 -24 1574 -16
rect -30 -33 665 -29
rect -30 -41 617 -37
rect 1522 -43 1526 -24
rect 1708 -43 1712 -24
rect -30 -49 569 -45
rect 1522 -47 1910 -43
rect -30 -57 139 -53
rect -30 -65 91 -61
rect -30 -73 43 -69
rect 11 -81 55 -77
rect 59 -81 103 -77
rect 107 -81 605 -77
rect 609 -81 653 -77
rect 657 -81 701 -77
rect 705 -81 1055 -77
rect 1059 -81 1103 -77
rect 1107 -81 1151 -77
rect 1155 -81 1917 -77
rect 146 -90 569 -85
rect 709 -90 1017 -85
rect 1160 -90 1345 -85
rect 1387 -90 1480 -85
rect 1574 -90 1667 -85
rect 1713 -90 1891 -85
<< polycontact >>
rect 334 525 338 529
<< m2contact >>
rect 1924 719 1933 724
rect 1162 707 1166 711
rect 1162 612 1166 616
rect 715 587 719 591
rect 460 529 464 533
rect 452 492 456 496
rect 460 493 464 497
rect 902 587 906 591
rect 715 493 719 497
rect 1162 587 1166 591
rect 1162 551 1166 555
rect 1891 659 1900 665
rect 1891 539 1900 545
rect 902 493 906 497
rect 910 529 914 533
rect 910 493 914 497
rect 1716 429 1720 433
rect 1723 411 1727 415
rect 1730 309 1734 313
rect 1737 291 1741 295
rect 1730 283 1734 287
rect 1723 261 1727 265
rect 1716 219 1720 223
rect 1716 77 1720 81
rect 1723 43 1727 47
rect 1737 197 1741 201
rect 1744 189 1748 193
rect 1751 459 1755 463
rect 1924 599 1933 605
rect 1891 419 1900 425
rect 1751 171 1755 175
rect 1758 381 1762 385
rect 1737 99 1741 103
rect 1758 69 1762 73
rect 1765 339 1769 343
rect 1761 51 1765 55
rect 1891 299 1900 305
rect 1891 179 1900 185
rect 1891 59 1900 65
rect 1730 21 1734 25
rect 342 0 346 4
rect 816 0 820 4
rect 1266 0 1270 4
rect 1067 -17 1071 -13
rect 1115 -18 1119 -14
rect 1019 -25 1023 -21
rect 665 -33 669 -29
rect 617 -41 621 -37
rect 569 -49 573 -45
rect 139 -57 143 -53
rect 91 -65 95 -61
rect 43 -73 47 -69
rect 7 -81 11 -77
rect 55 -81 59 -77
rect 103 -81 107 -77
rect 605 -81 609 -77
rect 653 -81 657 -77
rect 701 -81 705 -77
rect 1055 -81 1059 -77
rect 1103 -81 1107 -77
rect 1151 -81 1155 -77
rect 1903 -16 1907 -12
rect 1910 -47 1914 -43
rect 1924 479 1933 484
rect 1924 359 1933 365
rect 1924 239 1933 245
rect 1924 119 1933 125
rect 1924 0 1933 5
rect 1917 -81 1921 -77
rect 1891 -90 1900 -85
use IObuffertile IObuffertile_0
timestamp 951457029
transform 1 0 -67 0 1 -26
box 35 26 68 510
use pp1 pp1_0
timestamp 951985653
transform 1 0 0 0 1 0
box 0 0 441 544
use pp2 pp2_0
timestamp 951985653
transform 1 0 444 0 1 0
box -3 0 446 604
use pp3 pp3_0
timestamp 951985653
transform 1 0 894 0 1 0
box -3 0 446 724
use clockqual clockqual_0
timestamp 951296688
transform 1 0 -103 0 1 -35
box 103 -55 154 39
use clockqual clockqual_1
timestamp 951296688
transform 1 0 -55 0 1 -35
box 103 -55 154 39
use clockqual clockqual_2
timestamp 951296688
transform 1 0 -7 0 1 -35
box 103 -55 154 39
use clockqual clockqual_5
timestamp 951296688
transform -1 0 719 0 1 -35
box 103 -55 154 39
use clockqual clockqual_4
timestamp 951296688
transform -1 0 767 0 1 -35
box 103 -55 154 39
use clockqual clockqual_3
timestamp 951296688
transform -1 0 815 0 1 -35
box 103 -55 154 39
use clockqual clockqual_6
timestamp 951296688
transform -1 0 1169 0 1 -35
box 103 -55 154 39
use clockqual clockqual_7
timestamp 951296688
transform -1 0 1217 0 1 -35
box 103 -55 154 39
use clockqual clockqual_8
timestamp 951296688
transform -1 0 1265 0 1 -35
box 103 -55 154 39
use totalSR totalSR_0
timestamp 951985653
transform 1 0 1340 0 1 0
box 0 -8 375 724
use fullendmux fullendmux_0
timestamp 951985653
transform 1 0 1769 0 1 0
box 0 0 90 484
use IObuffertile IObuffertile_1
timestamp 951457029
transform 1 0 1821 0 1 -26
box 35 26 68 510
use SRclkdriver SRclkdriver_0
timestamp 951289694
transform 1 0 1340 0 1 -10
box 0 -80 51 14
use SRclkdriver SRclkdriver_1
timestamp 951289694
transform 1 0 1478 0 1 -10
box 0 -80 51 14
use SRclkdriver SRclkdriver_2
timestamp 951289694
transform 1 0 1526 0 1 -10
box 0 -80 51 14
use SRclkdriver SRclkdriver_3
timestamp 951289694
transform 1 0 1664 0 1 -10
box 0 -80 51 14
<< labels >>
rlabel metal2 1530 679 1530 679 3 SR_toControl_s1[19]
rlabel metal2 1530 645 1530 645 3 SR_toControl_s1[18]
rlabel metal2 1530 559 1530 559 3 SR_toControl_s1[17]
rlabel metal2 1530 525 1530 525 3 SR_toControl_s1[16]
rlabel metal1 1718 486 1718 486 7 SR_toControl_s1[15]
rlabel metal1 1725 486 1725 486 8 SR_toControl_s1[14]
rlabel metal1 1732 486 1732 486 1 SR_toControl_s1[13]
rlabel metal1 1739 486 1739 486 2 SR_toControl_s1[12]
rlabel metal1 1746 486 1746 486 3 SR_toControl_s1[11]
rlabel metal1 336 545 336 545 1 No_Connect_0
rlabel metal1 817 606 817 606 1 No_Connect_1
rlabel metal1 1267 726 1267 726 1 No_Connect_2
rlabel metal1 997 486 997 486 1 Kernel_Mux_s1[0]
rlabel metal1 961 486 961 486 3 Kernel_Mux_s1[1]
rlabel metal1 954 486 954 486 7 Kernel_Mux_s1[2]
rlabel metal1 1411 725 1411 725 1 Shift_Right_s2
rlabel metal1 1447 725 1447 725 8 Reset_Shift_s2
rlabel metal1 1454 725 1454 725 2 No_Shift_s2
rlabel metal1 266 503 266 503 8 pixel_bit0_v1
rlabel metal1 446 505 446 505 2 pixel_bit1_v1
rlabel metal1 896 506 896 506 2 pixel_bit2_v1
rlabel metal1 1832 485 1832 485 3 Sat_Control_s1[0]
rlabel metal1 1789 485 1789 485 8 Sat_Control_s1[1]
rlabel metal1 1825 485 1825 485 8 Sat_Control_s1[2]
rlabel metal1 1929 177 1929 177 3 Gnd
rlabel metal1 1895 165 1895 165 3 Vdd
rlabel metal1 1912 474 1912 474 1 Phi2
rlabel metal1 1904 467 1904 467 1 Phi1
rlabel metal1 1919 477 1919 477 4 Kernel_en_s1
rlabel metal2 1895 22 1895 22 3 Final_Output_s1[0]
rlabel metal2 1895 102 1895 102 3 Final_Output_s1[1]
rlabel metal2 1895 142 1895 142 3 Final_Output_s1[2]
rlabel metal2 1894 222 1894 222 3 Final_Output_s1[3]
rlabel metal2 1895 262 1895 262 3 Final_Output_s1[4]
rlabel metal2 1895 342 1895 342 3 Final_Output_s1[5]
rlabel metal2 1895 382 1895 382 3 Final_Output_s1[6]
rlabel metal2 1895 462 1895 462 3 Final_Output_s1[7]
rlabel metal2 -28 -71 -28 -71 7 Word_line_q1[0]
rlabel metal2 -28 -63 -28 -63 7 Word_line_q1[1]
rlabel metal2 -28 -55 -28 -55 7 Word_line_q1[2]
rlabel metal2 -28 -47 -28 -47 7 Word_line_q1[5]
rlabel metal2 -28 -39 -28 -39 7 Word_line_q1[4]
rlabel metal2 -28 -31 -28 -31 7 Word_line_q1[3]
rlabel metal2 -28 -23 -28 -23 7 Word_line_q1[8]
rlabel metal2 -28 -15 -28 -15 7 Word_line_q1[7]
rlabel metal2 -28 -7 -28 -7 7 Word_line_q1[6]
rlabel metal2 -31 24 -31 24 7 Kernel_Bus_b_v1[0]
rlabel metal2 -31 460 -31 460 7 Kernel_Bus_b_v1[7]
rlabel metal2 -31 384 -31 384 7 Kernel_Bus_b_v1[6]
rlabel metal2 -32 340 -32 340 7 Kernel_Bus_b_v1[5]
rlabel metal2 -31 264 -31 264 7 Kernel_Bus_b_v1[4]
rlabel metal2 -32 220 -32 220 7 Kernel_Bus_b_v1[3]
rlabel metal2 -32 144 -32 144 7 Kernel_Bus_b_v1[2]
rlabel metal2 -33 100 -33 100 7 Kernel_Bus_b_v1[1]
<< end >>
