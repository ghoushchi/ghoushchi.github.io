magic
tech scmos
timestamp 950486748
<< polysilicon >>
rect 71 114 86 150
rect 33 100 125 114
rect 71 62 86 100
<< metal1 >>
rect 0 167 168 335
rect 204 130 327 131
rect 204 126 312 130
rect 316 126 317 130
rect 321 126 322 130
rect 326 126 327 130
rect 204 125 327 126
rect 204 121 312 125
rect 316 121 317 125
rect 321 121 322 125
rect 326 121 327 125
rect 204 120 327 121
rect 204 116 312 120
rect 316 116 317 120
rect 321 116 322 120
rect 326 116 327 120
rect 204 115 327 116
rect 204 111 312 115
rect 316 111 317 115
rect 321 111 322 115
rect 326 111 327 115
rect 204 110 327 111
rect 204 106 312 110
rect 316 106 317 110
rect 321 106 322 110
rect 326 106 327 110
rect 204 105 327 106
rect 204 101 312 105
rect 316 101 317 105
rect 321 101 322 105
rect 326 101 327 105
rect 204 100 327 101
rect 204 96 312 100
rect 316 96 317 100
rect 321 96 322 100
rect 326 96 327 100
rect 204 95 327 96
rect 204 91 312 95
rect 316 91 317 95
rect 321 91 322 95
rect 326 91 327 95
rect 204 90 327 91
rect 204 86 312 90
rect 316 86 317 90
rect 321 86 322 90
rect 326 86 327 90
rect 204 85 327 86
rect 204 79 323 85
rect 204 13 254 79
rect 204 9 205 13
rect 209 9 210 13
rect 214 9 215 13
rect 219 9 220 13
rect 224 9 225 13
rect 229 9 230 13
rect 234 9 235 13
rect 239 9 240 13
rect 244 9 245 13
rect 249 9 254 13
rect 204 8 254 9
rect 204 4 205 8
rect 209 4 210 8
rect 214 4 215 8
rect 219 4 220 8
rect 224 4 225 8
rect 229 4 230 8
rect 234 4 235 8
rect 239 4 240 8
rect 244 4 245 8
rect 249 7 254 8
rect 272 55 308 59
rect 272 54 299 55
rect 272 46 289 54
rect 272 42 276 46
rect 280 42 281 46
rect 285 42 289 46
rect 272 41 289 42
rect 272 37 276 41
rect 280 37 281 41
rect 285 37 289 41
rect 272 10 289 37
rect 297 47 299 54
rect 307 47 308 55
rect 297 10 308 47
rect 272 7 308 10
rect 314 21 321 79
rect 314 20 323 21
rect 314 16 315 20
rect 314 15 319 16
rect 314 7 315 15
rect 249 4 250 7
<< metal2 >>
rect 1 330 303 334
rect 1 172 5 330
rect 163 172 303 330
rect 1 168 303 172
rect 167 73 303 168
rect 312 130 330 131
rect 316 126 317 130
rect 321 126 322 130
rect 326 126 330 130
rect 312 125 330 126
rect 316 121 317 125
rect 321 121 322 125
rect 326 121 330 125
rect 312 120 330 121
rect 316 116 317 120
rect 321 116 322 120
rect 326 116 330 120
rect 312 115 330 116
rect 316 111 317 115
rect 321 111 322 115
rect 326 111 330 115
rect 312 110 330 111
rect 316 106 317 110
rect 321 106 322 110
rect 326 106 330 110
rect 312 105 330 106
rect 316 101 317 105
rect 321 101 322 105
rect 326 101 330 105
rect 312 100 330 101
rect 316 96 317 100
rect 321 96 322 100
rect 326 96 330 100
rect 312 95 330 96
rect 316 91 317 95
rect 321 91 322 95
rect 326 91 330 95
rect 312 90 330 91
rect 316 86 317 90
rect 321 86 322 90
rect 326 86 330 90
rect 312 85 330 86
rect 167 46 330 73
rect 167 42 276 46
rect 280 42 281 46
rect 285 42 330 46
rect 167 41 330 42
rect 167 37 276 41
rect 280 37 281 41
rect 285 37 330 41
rect 167 25 330 37
rect 167 22 310 25
rect 204 9 205 13
rect 209 9 210 13
rect 214 9 215 13
rect 219 9 220 13
rect 224 9 225 13
rect 229 9 230 13
rect 234 9 235 13
rect 239 9 240 13
rect 244 9 245 13
rect 249 9 250 13
rect 204 8 250 9
rect 204 4 205 8
rect 209 4 210 8
rect 214 4 215 8
rect 219 4 220 8
rect 224 4 225 8
rect 229 4 230 8
rect 234 4 235 8
rect 239 4 240 8
rect 244 4 245 8
rect 249 4 250 8
rect 204 0 250 4
rect 262 0 310 22
rect 314 20 330 21
rect 314 16 315 20
rect 319 16 323 20
rect 327 16 330 20
rect 314 15 330 16
rect 314 11 320 15
rect 314 7 315 11
rect 319 7 320 11
rect 314 0 320 7
<< m2contact >>
rect 312 126 316 130
rect 317 126 321 130
rect 322 126 326 130
rect 312 121 316 125
rect 317 121 321 125
rect 322 121 326 125
rect 312 116 316 120
rect 317 116 321 120
rect 322 116 326 120
rect 312 111 316 115
rect 317 111 321 115
rect 322 111 326 115
rect 312 106 316 110
rect 317 106 321 110
rect 322 106 326 110
rect 312 101 316 105
rect 317 101 321 105
rect 322 101 326 105
rect 312 96 316 100
rect 317 96 321 100
rect 322 96 326 100
rect 312 91 316 95
rect 317 91 321 95
rect 322 91 326 95
rect 312 86 316 90
rect 317 86 321 90
rect 322 86 326 90
rect 205 9 209 13
rect 210 9 214 13
rect 215 9 219 13
rect 220 9 224 13
rect 225 9 229 13
rect 230 9 234 13
rect 235 9 239 13
rect 240 9 244 13
rect 245 9 249 13
rect 205 4 209 8
rect 210 4 214 8
rect 215 4 219 8
rect 220 4 224 8
rect 225 4 229 8
rect 230 4 234 8
rect 235 4 239 8
rect 240 4 244 8
rect 245 4 249 8
rect 276 42 280 46
rect 281 42 285 46
rect 276 37 280 41
rect 281 37 285 41
rect 315 16 319 20
rect 323 16 327 20
rect 315 7 319 11
<< psubstratepcontact >>
rect 319 16 323 20
rect 315 11 319 15
<< nsubstratencontact >>
rect 289 10 297 54
rect 299 47 307 55
<< psubstratepdiff >>
rect 314 20 330 21
rect 314 16 319 20
rect 323 16 330 20
rect 314 15 330 16
rect 314 11 315 15
rect 319 11 320 15
rect 314 0 320 11
<< nsubstratendiff >>
rect 264 55 330 71
rect 264 54 299 55
rect 264 10 289 54
rect 297 47 299 54
rect 307 47 330 55
rect 297 27 330 47
rect 297 10 308 27
rect 264 0 308 10
<< pad >>
rect 5 172 163 330
<< glass >>
rect 11 178 157 324
<< labels >>
rlabel metal2 286 57 286 57 6 Vdd
rlabel metal1 0 335 0 335 4 sllu
rlabel space 0 0 0 0 2 sllu_1988
rlabel space 330 335 330 335 6 sllu_1988
rlabel metal2 330 73 330 73 6 {e}tiny12_b
rlabel metal2 330 85 330 85 6 {e}tiny12_t
rlabel metal2 250 0 250 0 8 {s}tiny12_t
rlabel metal2 262 0 262 0 8 {s}tiny12_b
rlabel metal2 330 115 330 115 6 {e}*
rlabel metal2 220 0 220 0 8 {s}*
<< end >>
