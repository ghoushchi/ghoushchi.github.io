magic
tech scmos
timestamp 950486748
<< metal1 >>
rect 67 168 219 320
rect 11 101 12 105
rect 260 101 261 105
rect 18 50 262 58
rect 18 46 20 50
rect 24 46 25 50
rect 29 46 30 50
rect 34 46 35 50
rect 39 48 262 50
rect 39 46 237 48
rect 18 45 237 46
rect 18 41 20 45
rect 24 41 25 45
rect 29 41 30 45
rect 34 41 35 45
rect 39 44 237 45
rect 241 44 242 48
rect 246 44 247 48
rect 251 44 252 48
rect 256 44 257 48
rect 261 44 262 48
rect 39 43 262 44
rect 39 41 237 43
rect 18 40 237 41
rect 18 36 20 40
rect 24 36 25 40
rect 29 36 30 40
rect 34 36 35 40
rect 39 39 237 40
rect 241 39 242 43
rect 246 39 247 43
rect 251 39 252 43
rect 256 39 257 43
rect 261 39 262 43
rect 39 38 262 39
rect 39 36 237 38
rect 18 35 237 36
rect 18 31 20 35
rect 24 31 25 35
rect 29 31 30 35
rect 34 31 35 35
rect 39 34 237 35
rect 241 34 242 38
rect 246 34 247 38
rect 251 34 252 38
rect 256 34 257 38
rect 261 34 262 38
rect 39 33 262 34
rect 39 31 237 33
rect 18 30 237 31
rect 18 26 20 30
rect 24 26 25 30
rect 29 26 30 30
rect 34 26 35 30
rect 39 29 237 30
rect 241 29 242 33
rect 246 29 247 33
rect 251 29 252 33
rect 256 29 257 33
rect 261 29 262 33
rect 39 28 262 29
rect 39 26 237 28
rect 18 25 237 26
rect 18 21 20 25
rect 24 21 25 25
rect 29 21 30 25
rect 34 21 35 25
rect 39 24 237 25
rect 241 24 242 28
rect 246 24 247 28
rect 251 24 252 28
rect 256 24 257 28
rect 261 24 262 28
rect 39 23 262 24
rect 39 21 237 23
rect 18 19 237 21
rect 241 19 242 23
rect 246 19 247 23
rect 251 19 252 23
rect 256 19 257 23
rect 261 19 262 23
rect 18 17 262 19
rect 258 13 262 17
rect 18 10 262 13
rect 41 5 240 6
rect 68 1 72 5
rect 76 1 80 5
rect 84 1 88 5
rect 92 1 96 5
rect 100 1 104 5
rect 108 1 112 5
rect 116 1 120 5
rect 124 1 128 5
rect 132 1 136 5
rect 140 1 144 5
rect 148 1 152 5
rect 156 1 160 5
rect 164 1 168 5
rect 172 1 176 5
rect 180 1 184 5
rect 188 1 192 5
rect 196 1 200 5
rect 204 1 208 5
rect 212 1 216 5
rect 220 1 224 5
rect 41 0 240 1
<< metal2 >>
rect 68 315 218 319
rect 68 173 72 315
rect 214 173 218 315
rect 68 169 218 173
rect 68 116 219 169
rect 0 70 285 116
rect 0 50 39 58
rect 0 46 20 50
rect 24 46 25 50
rect 29 46 30 50
rect 34 46 35 50
rect 0 45 39 46
rect 0 41 20 45
rect 24 41 25 45
rect 29 41 30 45
rect 34 41 35 45
rect 0 40 39 41
rect 0 36 20 40
rect 24 36 25 40
rect 29 36 30 40
rect 34 36 35 40
rect 0 35 39 36
rect 0 31 20 35
rect 24 31 25 35
rect 29 31 30 35
rect 34 31 35 35
rect 0 30 39 31
rect 0 26 20 30
rect 24 26 25 30
rect 29 26 30 30
rect 34 26 35 30
rect 0 25 39 26
rect 0 21 20 25
rect 24 21 25 25
rect 29 21 30 25
rect 34 21 35 25
rect 0 10 39 21
rect 68 6 219 70
rect 237 48 285 58
rect 241 44 242 48
rect 246 44 247 48
rect 251 44 252 48
rect 256 44 257 48
rect 261 44 285 48
rect 237 43 285 44
rect 241 39 242 43
rect 246 39 247 43
rect 251 39 252 43
rect 256 39 257 43
rect 261 39 285 43
rect 237 38 285 39
rect 241 34 242 38
rect 246 34 247 38
rect 251 34 252 38
rect 256 34 257 38
rect 261 34 285 38
rect 237 33 285 34
rect 241 29 242 33
rect 246 29 247 33
rect 251 29 252 33
rect 256 29 257 33
rect 261 29 285 33
rect 237 28 285 29
rect 241 24 242 28
rect 246 24 247 28
rect 251 24 252 28
rect 256 24 257 28
rect 261 24 285 28
rect 237 23 285 24
rect 241 19 242 23
rect 246 19 247 23
rect 251 19 252 23
rect 256 19 257 23
rect 261 19 285 23
rect 237 10 285 19
rect 0 5 285 6
rect 0 1 40 5
rect 44 1 48 5
rect 52 1 56 5
rect 60 1 228 5
rect 232 1 236 5
rect 240 1 244 5
rect 248 1 252 5
rect 256 1 260 5
rect 264 1 268 5
rect 272 1 285 5
rect 0 0 285 1
<< m2contact >>
rect 20 46 24 50
rect 25 46 29 50
rect 30 46 34 50
rect 35 46 39 50
rect 20 41 24 45
rect 25 41 29 45
rect 30 41 34 45
rect 35 41 39 45
rect 237 44 241 48
rect 242 44 246 48
rect 247 44 251 48
rect 252 44 256 48
rect 257 44 261 48
rect 20 36 24 40
rect 25 36 29 40
rect 30 36 34 40
rect 35 36 39 40
rect 237 39 241 43
rect 242 39 246 43
rect 247 39 251 43
rect 252 39 256 43
rect 257 39 261 43
rect 20 31 24 35
rect 25 31 29 35
rect 30 31 34 35
rect 35 31 39 35
rect 237 34 241 38
rect 242 34 246 38
rect 247 34 251 38
rect 252 34 256 38
rect 257 34 261 38
rect 20 26 24 30
rect 25 26 29 30
rect 30 26 34 30
rect 35 26 39 30
rect 237 29 241 33
rect 242 29 246 33
rect 247 29 251 33
rect 252 29 256 33
rect 257 29 261 33
rect 20 21 24 25
rect 25 21 29 25
rect 30 21 34 25
rect 35 21 39 25
rect 237 24 241 28
rect 242 24 246 28
rect 247 24 251 28
rect 252 24 256 28
rect 257 24 261 28
rect 237 19 241 23
rect 242 19 246 23
rect 247 19 251 23
rect 252 19 256 23
rect 257 19 261 23
rect 40 1 44 5
rect 48 1 52 5
rect 56 1 60 5
rect 228 1 232 5
rect 236 1 240 5
rect 244 1 248 5
rect 252 1 256 5
rect 260 1 264 5
rect 268 1 272 5
<< psubstratepcontact >>
rect 12 101 260 105
rect 44 1 48 5
rect 52 1 56 5
rect 60 1 68 5
rect 72 1 76 5
rect 80 1 84 5
rect 88 1 92 5
rect 96 1 100 5
rect 104 1 108 5
rect 112 1 116 5
rect 120 1 124 5
rect 128 1 132 5
rect 136 1 140 5
rect 144 1 148 5
rect 152 1 156 5
rect 160 1 164 5
rect 168 1 172 5
rect 176 1 180 5
rect 184 1 188 5
rect 192 1 196 5
rect 200 1 204 5
rect 208 1 212 5
rect 216 1 220 5
rect 224 1 228 5
rect 232 1 236 5
rect 240 1 244 5
rect 248 1 252 5
rect 256 1 260 5
rect 264 1 268 5
rect 272 1 276 5
<< nsubstratencontact >>
rect 18 13 258 17
<< psubstratepdiff >>
rect 4 139 281 141
rect 0 133 285 139
rect 0 105 8 133
rect 131 107 160 133
rect 254 107 285 133
rect 131 105 285 107
rect 0 101 12 105
rect 260 101 285 105
rect 0 100 285 101
rect 43 80 47 100
rect 67 80 74 100
rect 187 80 195 100
rect 43 76 195 80
rect 0 5 285 6
rect 0 1 44 5
rect 48 1 52 5
rect 56 1 60 5
rect 68 1 72 5
rect 76 1 80 5
rect 84 1 88 5
rect 92 1 96 5
rect 100 1 104 5
rect 108 1 112 5
rect 116 1 120 5
rect 124 1 128 5
rect 132 1 136 5
rect 140 1 144 5
rect 148 1 152 5
rect 156 1 160 5
rect 164 1 168 5
rect 172 1 176 5
rect 180 1 184 5
rect 188 1 192 5
rect 196 1 200 5
rect 204 1 208 5
rect 212 1 216 5
rect 220 1 224 5
rect 228 1 232 5
rect 236 1 240 5
rect 244 1 248 5
rect 252 1 256 5
rect 260 1 264 5
rect 268 1 272 5
rect 276 1 285 5
rect 0 0 285 1
<< nsubstratendiff >>
rect 0 52 285 56
rect 0 46 6 52
rect 0 18 7 46
rect 43 18 47 52
rect 67 20 80 52
rect 131 50 141 52
rect 174 51 285 52
rect 174 20 188 51
rect 67 18 188 20
rect 272 18 285 51
rect 0 17 285 18
rect 0 13 18 17
rect 258 13 285 17
rect 0 12 285 13
<< pad >>
rect 72 173 214 315
<< glass >>
rect 78 179 208 309
<< labels >>
rlabel space 0 320 0 320 4 sllu_1988
rlabel space 285 320 285 320 6 mosis_tinychip
rlabel metal1 143 234 143 234 6 pad
rlabel metal2 0 70 0 70 4 {w}tiny12_t
rlabel metal2 0 58 0 58 4 {w}tiny12_b
rlabel metal2 285 70 285 70 6 {e}tiny12_t
rlabel metal2 285 58 285 58 6 {e}tiny12_b
rlabel metal2 143 0 143 0 8 .GND
rlabel psubstratepdiff 0 100 0 100 4 {w}*
rlabel psubstratepdiff 285 100 285 100 6 {e}*
<< end >>
