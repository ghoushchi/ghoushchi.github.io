magic
tech scmos
timestamp 951727448
<< m2contact >>
rect -2 -2 2 2
<< end >>
