magic
tech scmos
timestamp 830644267
<< pad >>
rect 5 3072 163 3230
rect 402 3088 544 3230
rect 686 3088 828 3230
rect 972 3088 1114 3230
rect 1256 3088 1398 3230
rect 1542 3088 1684 3230
rect 1826 3088 1968 3230
rect 2112 3088 2254 3230
rect 2396 3088 2538 3230
rect 2682 3088 2824 3230
rect 3062 3072 3220 3230
rect 5 2687 147 2829
rect 3078 2687 3220 2829
rect 5 2401 147 2543
rect 3078 2401 3220 2543
rect 5 2117 147 2259
rect 3078 2117 3220 2259
rect 5 1831 147 1973
rect 3078 1831 3220 1973
rect 5 1547 147 1689
rect 3078 1547 3220 1689
rect 5 1261 147 1403
rect 3078 1261 3220 1403
rect 5 977 147 1119
rect 3078 977 3220 1119
rect 5 691 147 833
rect 3078 691 3220 833
rect 5 407 147 549
rect 3078 407 3220 549
rect 5 5 163 163
rect 402 5 544 147
rect 686 5 828 147
rect 972 5 1114 147
rect 1256 5 1398 147
rect 1542 5 1684 147
rect 1826 5 1968 147
rect 2112 5 2254 147
rect 2396 5 2538 147
rect 2682 5 2824 147
rect 3062 5 3220 163
use chip chip_0
timestamp 789595518
transform 1 0 0 0 1 0
box 0 0 3225 3235
<< labels >>
rlabel pad 3062 3072 3220 3230 1 Pin5
rlabel pad 3078 2687 3220 2829 1 Pin4
rlabel pad 3078 2401 3220 2543 1 Pin3
rlabel pad 3078 2117 3220 2259 1 Pin2
rlabel pad 3078 1831 3220 1973 1 Pin1
rlabel pad 3078 1547 3220 1689 1 Pin40
rlabel pad 3078 1261 3220 1403 1 Pin39
rlabel pad 3078 977 3220 1119 1 Pin38
rlabel pad 3078 691 3220 833 1 Pin37
rlabel pad 3078 407 3220 549 1 Pin36
rlabel pad 3062 5 3220 163 1 Pin35
rlabel pad 2682 5 2824 147 1 Pin34
rlabel pad 2396 5 2538 147 1 Pin33
rlabel pad 2112 5 2254 147 1 Pin32
rlabel pad 1826 5 1968 147 1 Pin31
rlabel pad 1542 5 1684 147 1 Pin30
rlabel pad 1256 5 1398 147 1 Pin29
rlabel pad 972 5 1114 147 1 Pin28
rlabel pad 686 5 828 147 1 Pin27
rlabel pad 402 5 544 147 1 Pin26
rlabel pad 5 5 163 163 1 Pin25
rlabel pad 5 407 147 549 1 Pin24
rlabel pad 5 691 147 833 1 Pin23
rlabel pad 5 977 147 1119 1 Pin22
rlabel pad 5 1261 147 1403 1 Pin21
rlabel pad 5 1547 147 1689 1 Pin20
rlabel pad 5 1831 147 1973 1 Pin19
rlabel pad 5 2117 147 2259 1 Pin18
rlabel pad 5 2401 147 2543 1 Pin17
rlabel pad 5 2687 147 2829 1 Pin16
rlabel pad 5 3072 163 3230 1 Pin15
rlabel pad 402 3088 544 3230 1 Pin14
rlabel pad 686 3088 828 3230 1 Pin13
rlabel pad 972 3088 1114 3230 1 Pin12
rlabel pad 1256 3088 1398 3230 1 Pin11
rlabel pad 1542 3088 1684 3230 1 Pin10
rlabel pad 1826 3088 1968 3230 1 Pin9
rlabel pad 2112 3088 2254 3230 1 Pin8
rlabel pad 2396 3088 2538 3230 1 Pin7
rlabel pad 2682 3088 2824 3230 1 Pin6
<< end >>
