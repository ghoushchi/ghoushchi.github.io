magic
tech scmos
timestamp 950486748
use tl 2_0
timestamp 950486748
transform 1 0 0 0 1 2900
box 0 0 330 335
use io 3_0
timestamp 950486748
transform 1 0 330 0 1 2915
box 0 0 285 320
use io 3_1
timestamp 950486748
transform -1 0 900 0 1 2915
box 0 0 285 320
use io 3_2
timestamp 950486748
transform 1 0 900 0 1 2915
box 0 0 285 320
use io 3_3
timestamp 950486748
transform -1 0 1470 0 1 2915
box 0 0 285 320
use gnd 4_0
timestamp 950486748
transform 1 0 1470 0 1 2915
box 0 0 285 320
use io 3_4
timestamp 950486748
transform -1 0 2040 0 1 2915
box 0 0 285 320
use io 3_5
timestamp 950486748
transform 1 0 2040 0 1 2915
box 0 0 285 320
use io 3_6
timestamp 950486748
transform -1 0 2610 0 1 2915
box 0 0 285 320
use io 3_7
timestamp 950486748
transform 1 0 2610 0 1 2915
box 0 0 285 320
use tr 5_0
timestamp 950486748
transform 1 0 2895 0 1 2900
box 0 0 330 335
use io 3_8
timestamp 950486748
transform 0 -1 320 1 0 2615
box 0 0 285 320
use io 3_9
timestamp 950486748
transform 0 -1 320 -1 0 2615
box 0 0 285 320
use io 3_10
timestamp 950486748
transform 0 -1 320 1 0 2045
box 0 0 285 320
use io 3_11
timestamp 950486748
transform 0 -1 320 -1 0 2045
box 0 0 285 320
use io 3_12
timestamp 950486748
transform 0 -1 320 1 0 1475
box 0 0 285 320
use io 3_13
timestamp 950486748
transform 0 -1 320 -1 0 1475
box 0 0 285 320
use io 3_14
timestamp 950486748
transform 0 -1 320 1 0 905
box 0 0 285 320
use io 3_15
timestamp 950486748
transform 0 -1 320 -1 0 905
box 0 0 285 320
use io 3_16
timestamp 950486748
transform 0 -1 320 1 0 335
box 0 0 285 320
use io 3_17
timestamp 950486748
transform 0 1 2905 1 0 2615
box 0 0 285 320
use io 3_18
timestamp 950486748
transform 0 1 2905 -1 0 2615
box 0 0 285 320
use io 3_19
timestamp 950486748
transform 0 1 2905 1 0 2045
box 0 0 285 320
use io 3_20
timestamp 950486748
transform 0 1 2905 -1 0 2045
box 0 0 285 320
use io 3_21
timestamp 950486748
transform 0 1 2905 1 0 1475
box 0 0 285 320
use io 3_22
timestamp 950486748
transform 0 1 2905 -1 0 1475
box 0 0 285 320
use io 3_23
timestamp 950486748
transform 0 1 2905 1 0 905
box 0 0 285 320
use io 3_24
timestamp 950486748
transform 0 1 2905 -1 0 905
box 0 0 285 320
use io 3_25
timestamp 950486748
transform 0 1 2905 1 0 335
box 0 0 285 320
use bl 6_0
timestamp 950486748
transform 1 0 0 0 1 0
box 0 0 330 335
use io 3_26
timestamp 950486748
transform 1 0 330 0 -1 320
box 0 0 285 320
use io 3_27
timestamp 950486748
transform -1 0 900 0 -1 320
box 0 0 285 320
use io 3_28
timestamp 950486748
transform 1 0 900 0 -1 320
box 0 0 285 320
use io 3_29
timestamp 950486748
transform -1 0 1470 0 -1 320
box 0 0 285 320
use vdd 7_0
timestamp 950486748
transform 1 0 1470 0 -1 320
box 0 0 285 320
use io 3_30
timestamp 950486748
transform -1 0 2040 0 -1 320
box 0 0 285 320
use io 3_31
timestamp 950486748
transform 1 0 2040 0 -1 320
box 0 0 285 320
use io 3_32
timestamp 950486748
transform -1 0 2610 0 -1 320
box 0 0 285 320
use io 3_33
timestamp 950486748
transform 1 0 2610 0 -1 320
box 0 0 285 320
use br 8_0
timestamp 950486748
transform 1 0 2895 0 1 0
box 0 0 330 335
<< end >>
