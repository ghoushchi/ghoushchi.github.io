magic
tech scmos
timestamp 951727448
<< pwell >>
rect 0 0 48 32
<< nwell >>
rect 0 32 48 64
<< polysilicon >>
rect 11 52 13 54
rect 19 52 21 54
rect 27 52 29 54
rect 11 22 13 40
rect 15 22 17 24
rect 19 22 21 40
rect 27 39 29 40
rect 27 37 38 39
rect 25 27 29 29
rect 27 22 29 27
rect 31 22 33 37
rect 35 22 37 24
rect 11 6 13 14
rect 15 10 17 14
rect 19 12 21 14
rect 27 12 29 14
rect 31 10 33 14
rect 15 8 33 10
rect 35 6 37 14
rect 11 4 37 6
<< ndiffusion >>
rect 10 14 11 22
rect 13 14 15 22
rect 17 14 19 22
rect 21 14 22 22
rect 26 14 27 22
rect 29 14 31 22
rect 33 14 35 22
rect 37 14 38 22
<< pdiffusion >>
rect 10 40 11 52
rect 13 40 14 52
rect 18 40 19 52
rect 21 40 22 52
rect 26 40 27 52
rect 29 40 30 52
<< metal1 >>
rect 0 56 6 60
rect 10 56 22 60
rect 26 56 38 60
rect 42 56 48 60
rect 6 52 10 56
rect 22 52 26 56
rect 14 36 18 40
rect 7 31 10 32
rect 14 20 17 32
rect 22 31 25 32
rect 14 17 22 20
rect 30 20 33 40
rect 38 36 42 37
rect 26 17 33 20
rect 6 8 10 14
rect 38 8 42 14
rect 0 4 6 8
rect 10 4 38 8
rect 42 4 48 8
<< ntransistor >>
rect 11 14 13 22
rect 15 14 17 22
rect 19 14 21 22
rect 27 14 29 22
rect 31 14 33 22
rect 35 14 37 22
<< ptransistor >>
rect 11 40 13 52
rect 19 40 21 52
rect 27 40 29 52
<< polycontact >>
rect 7 27 11 31
rect 38 37 42 41
rect 21 27 25 31
<< ndcontact >>
rect 6 14 10 22
rect 22 14 26 22
rect 38 14 42 22
<< pdcontact >>
rect 6 40 10 52
rect 14 40 18 52
rect 22 40 26 52
rect 30 40 34 52
<< m2contact >>
rect 6 32 10 36
rect 14 32 18 36
rect 22 32 26 36
rect 38 32 42 36
<< psubstratepcontact >>
rect 6 4 10 8
rect 38 4 42 8
<< nsubstratencontact >>
rect 6 56 10 60
rect 22 56 26 60
rect 38 56 42 60
<< labels >>
rlabel m2contact 8 34 8 34 6 In2
rlabel m2contact 16 34 16 34 6 Out_b
rlabel m2contact 24 34 24 34 6 In0
rlabel metal1 4 6 4 6 6 GND
rlabel metal1 44 58 44 58 6 Vdd
rlabel metal1 4 58 4 58 6 Vdd
rlabel metal1 44 6 44 6 6 GND
rlabel m2contact 40 34 40 34 6 In1
<< end >>
