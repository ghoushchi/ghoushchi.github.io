magic
tech scmos
timestamp 951088720
<< nwell >>
rect 39 29 96 61
rect 40 20 96 29
<< polysilicon >>
rect 57 47 60 48
rect 53 46 60 47
rect 80 46 82 48
rect 55 42 60 44
rect 80 42 82 44
rect 55 28 57 42
rect 38 26 57 28
rect 64 26 67 28
rect 77 26 83 28
rect 55 18 57 26
rect 55 16 75 18
rect 53 12 67 13
rect 57 11 67 12
rect 65 10 67 11
rect 73 10 75 16
rect 81 10 83 26
rect 39 -3 41 5
rect 65 3 67 5
rect 73 3 75 5
rect 81 3 83 5
<< ndiffusion >>
rect 64 5 65 10
rect 67 5 68 10
rect 72 5 73 10
rect 75 5 76 10
rect 80 5 81 10
rect 83 5 84 10
<< pdiffusion >>
rect 60 48 80 49
rect 60 44 80 46
rect 60 41 80 42
rect 67 28 77 29
rect 67 25 77 26
<< metal1 >>
rect 39 34 43 61
rect 46 33 50 61
rect 53 51 57 61
rect 65 57 75 61
rect 60 53 80 57
rect 80 49 88 53
rect 46 29 47 33
rect 39 9 43 10
rect 46 -3 50 29
rect 54 12 57 47
rect 60 30 63 37
rect 84 33 88 49
rect 77 29 88 33
rect 60 17 63 26
rect 77 22 84 25
rect 60 14 72 17
rect 68 10 72 14
rect 84 10 88 21
rect 53 -3 56 8
rect 60 1 64 5
rect 76 1 80 5
rect 64 -3 65 1
rect 69 -3 80 1
<< metal2 >>
rect 39 57 75 61
rect 80 57 96 61
rect 39 56 96 57
rect -17 48 143 52
rect -17 38 143 42
rect 51 29 143 33
rect -17 22 36 26
rect 88 21 112 25
rect 140 22 143 29
rect 8 14 25 18
rect 21 10 39 14
rect 39 1 96 2
rect 39 -3 65 1
rect 69 -3 96 1
<< ntransistor >>
rect 65 5 67 10
rect 73 5 75 10
rect 81 5 83 10
<< ptransistor >>
rect 60 46 80 48
rect 60 42 80 44
rect 67 26 77 28
<< polycontact >>
rect 53 47 57 51
rect 34 25 38 29
rect 60 26 64 30
rect 39 5 43 9
rect 53 8 57 12
<< ndcontact >>
rect 60 5 64 10
rect 68 5 72 10
rect 76 5 80 10
rect 84 5 88 10
<< pdcontact >>
rect 60 49 80 53
rect 60 37 80 41
rect 67 29 77 33
rect 67 21 77 25
<< m2contact >>
rect 75 57 80 61
rect 47 29 51 33
rect 32 18 36 22
rect 4 14 8 18
rect 39 10 43 14
rect 84 21 88 25
rect 112 21 116 25
rect 140 18 144 22
rect 65 -3 69 1
<< psubstratepcontact >>
rect 60 -3 64 1
<< nsubstratencontact >>
rect 60 57 65 61
use InvLatch InvLatch_0
timestamp 951088720
transform 1 0 -11 0 1 -3
box -1 0 50 64
use InvLatch InvLatch_1
timestamp 951088720
transform 1 0 97 0 1 -3
box -1 0 50 64
<< labels >>
rlabel metal2 -15 50 -15 50 3 random1
rlabel metal2 -16 40 -16 40 3 random2
rlabel metal1 48 55 48 55 1 to_bottom
rlabel metal1 55 54 55 54 1 Set
rlabel metal2 80 -2 80 -2 1 Gnd
rlabel metal2 -15 24 -15 24 3 Output
rlabel metal2 92 59 92 59 5 Vdd
<< end >>
