magic
tech scmos
timestamp 950486748
<< polysilicon >>
rect 37 218 123 232
<< metal1 >>
rect 244 327 245 331
rect 249 328 250 331
rect 249 327 315 328
rect 240 326 315 327
rect 244 322 245 326
rect 249 324 315 326
rect 313 320 315 324
rect 313 319 319 320
rect 283 296 291 298
rect 280 292 281 296
rect 285 292 286 296
rect 290 294 291 296
rect 313 315 315 319
rect 290 293 303 294
rect 290 292 295 293
rect 276 291 295 292
rect 280 287 281 291
rect 285 287 286 291
rect 290 287 295 291
rect 276 286 295 287
rect 280 282 281 286
rect 285 282 286 286
rect 290 282 295 286
rect 313 250 323 315
rect 313 249 327 250
rect 317 245 318 249
rect 322 245 323 249
rect 313 244 327 245
rect 317 240 318 244
rect 322 240 323 244
rect 0 0 168 168
<< metal2 >>
rect 204 331 250 335
rect 204 327 240 331
rect 244 327 245 331
rect 249 327 250 331
rect 204 326 250 327
rect 204 322 240 326
rect 244 322 245 326
rect 249 322 250 326
rect 204 250 250 322
rect 262 310 310 335
rect 314 328 320 335
rect 314 324 315 328
rect 319 324 320 328
rect 314 320 320 324
rect 314 319 330 320
rect 314 315 315 319
rect 319 315 323 319
rect 327 315 330 319
rect 314 314 330 315
rect 262 296 330 310
rect 262 292 276 296
rect 280 292 281 296
rect 285 292 286 296
rect 290 292 330 296
rect 262 291 330 292
rect 262 287 276 291
rect 280 287 281 291
rect 285 287 286 291
rect 290 287 330 291
rect 262 286 330 287
rect 262 282 276 286
rect 280 282 281 286
rect 285 282 286 286
rect 290 282 330 286
rect 262 262 330 282
rect 204 249 330 250
rect 204 245 313 249
rect 317 245 318 249
rect 322 245 323 249
rect 327 245 330 249
rect 204 244 330 245
rect 204 240 313 244
rect 317 240 318 244
rect 322 240 323 244
rect 327 240 330 244
rect 204 204 330 240
rect 204 167 303 204
rect 1 163 303 167
rect 1 5 5 163
rect 163 5 303 163
rect 1 1 303 5
<< m2contact >>
rect 240 327 244 331
rect 245 327 249 331
rect 240 322 244 326
rect 245 322 249 326
rect 315 324 319 328
rect 276 292 280 296
rect 281 292 285 296
rect 286 292 290 296
rect 315 315 319 319
rect 323 315 327 319
rect 276 287 280 291
rect 281 287 285 291
rect 286 287 290 291
rect 276 282 280 286
rect 281 282 285 286
rect 286 282 290 286
rect 313 245 317 249
rect 318 245 322 249
rect 323 245 327 249
rect 313 240 317 244
rect 318 240 322 244
rect 323 240 327 244
<< psubstratepcontact >>
rect 315 320 319 324
rect 319 315 323 319
<< nsubstratencontact >>
rect 283 298 291 318
rect 295 277 303 293
<< psubstratepdiff >>
rect 314 324 320 335
rect 314 320 315 324
rect 319 320 320 324
rect 314 319 330 320
rect 314 315 319 319
rect 323 315 330 319
rect 314 314 330 315
<< nsubstratendiff >>
rect 268 318 302 335
rect 268 298 283 318
rect 291 303 302 318
rect 291 298 330 303
rect 268 293 330 298
rect 268 277 295 293
rect 303 277 330 293
rect 268 269 330 277
<< pad >>
rect 5 5 163 163
<< glass >>
rect 11 11 157 157
<< labels >>
rlabel metal2 286 278 286 278 6 Vdd
rlabel metal1 0 0 0 0 2 sllu
rlabel space 0 335 0 335 4 sllu_1988
rlabel space 330 0 330 0 8 sllu_1988
rlabel metal2 253 207 253 207 6 GND
rlabel space 90 263 90 263 6 Copy_Righted_MOSIS
rlabel space 90 253 90 253 6 Shih_Lien_Lu
rlabel space 90 245 90 245 6 1988
rlabel metal2 330 250 330 250 6 {e}tiny12_t
rlabel metal2 330 262 330 262 6 {e}tiny12_b
rlabel metal2 250 335 250 335 6 {n}tiny12_t
rlabel metal2 262 335 262 335 6 {n}tiny12_b
rlabel metal2 330 220 330 220 6 {e}*
rlabel metal2 204 335 204 335 6 {n}*
<< end >>
