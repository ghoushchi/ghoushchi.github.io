magic
tech scmos
timestamp 951963504
<< polysilicon >>
rect 0 -22 393 2
rect 0 -24 254 -22
rect 0 -26 18 -24
rect 33 -26 66 -24
rect 84 -26 121 -24
rect 133 -26 254 -24
rect 0 -32 16 -26
rect 37 -28 66 -26
rect 88 -28 117 -26
rect 20 -32 29 -30
rect 0 -38 31 -32
rect 39 -38 66 -28
rect 90 -30 115 -28
rect 0 -40 29 -38
rect 0 -44 27 -40
rect 37 -42 43 -38
rect 35 -44 43 -42
rect 57 -44 66 -38
rect 0 -46 23 -44
rect 33 -46 66 -44
rect 0 -48 20 -46
rect 31 -48 66 -46
rect 0 -50 18 -48
rect 29 -50 66 -48
rect 74 -32 82 -30
rect 74 -34 84 -32
rect 92 -34 113 -30
rect 123 -32 131 -30
rect 137 -32 254 -26
rect 121 -34 135 -32
rect 137 -34 148 -32
rect 160 -34 168 -32
rect 176 -34 180 -32
rect 188 -34 195 -32
rect 203 -34 213 -32
rect 221 -34 229 -32
rect 242 -34 254 -32
rect 74 -46 86 -34
rect 94 -46 111 -34
rect 119 -36 145 -34
rect 162 -36 168 -34
rect 191 -36 197 -34
rect 119 -38 143 -36
rect 164 -38 168 -36
rect 119 -46 141 -38
rect 152 -40 156 -38
rect 74 -48 84 -46
rect 74 -50 82 -48
rect 92 -50 113 -46
rect 121 -48 135 -46
rect 123 -50 131 -48
rect 137 -50 141 -46
rect 150 -48 158 -40
rect 152 -50 156 -48
rect 166 -50 168 -38
rect 0 -56 16 -50
rect 41 -56 66 -50
rect 90 -52 115 -50
rect 137 -52 143 -50
rect 164 -52 168 -50
rect 86 -54 117 -52
rect 137 -54 145 -52
rect 82 -56 121 -54
rect 133 -56 148 -54
rect 160 -56 168 -52
rect 176 -56 184 -38
rect 193 -40 197 -36
rect 205 -40 211 -34
rect 219 -36 227 -34
rect 244 -36 254 -34
rect 219 -38 225 -36
rect 246 -38 254 -36
rect 219 -40 223 -38
rect 234 -40 238 -38
rect 193 -46 199 -40
rect 207 -46 209 -40
rect 217 -46 223 -40
rect 193 -52 201 -46
rect 213 -48 223 -46
rect 231 -48 240 -40
rect 215 -50 223 -48
rect 234 -50 238 -48
rect 248 -50 254 -38
rect 213 -52 225 -50
rect 246 -52 254 -50
rect 193 -56 203 -52
rect 213 -54 227 -52
rect 213 -56 229 -54
rect 242 -56 254 -52
rect 262 -26 315 -22
rect 262 -32 295 -26
rect 303 -28 315 -26
rect 324 -28 393 -22
rect 303 -32 393 -28
rect 262 -52 264 -32
rect 272 -50 281 -32
rect 289 -38 293 -32
rect 309 -38 315 -32
rect 262 -54 266 -52
rect 289 -54 295 -38
rect 303 -50 315 -38
rect 262 -56 268 -54
rect 277 -56 281 -54
rect 289 -56 299 -54
rect 309 -56 315 -50
rect 324 -34 332 -32
rect 344 -34 354 -32
rect 363 -34 367 -32
rect 375 -34 393 -32
rect 324 -36 330 -34
rect 346 -36 354 -34
rect 377 -36 393 -34
rect 324 -38 328 -36
rect 348 -38 354 -36
rect 324 -50 326 -38
rect 336 -40 340 -38
rect 334 -48 342 -40
rect 336 -50 340 -48
rect 350 -50 354 -38
rect 324 -52 328 -50
rect 348 -52 354 -50
rect 324 -54 330 -52
rect 324 -56 332 -54
rect 344 -56 354 -52
rect 363 -56 371 -38
rect 379 -56 393 -36
rect 0 -75 393 -56
rect 0 -77 215 -75
rect 0 -110 129 -77
rect 152 -81 215 -77
rect 223 -81 393 -75
rect 152 -83 393 -81
rect 137 -85 393 -83
rect 137 -89 156 -85
rect 164 -87 168 -85
rect 176 -87 191 -85
rect 178 -89 188 -87
rect 150 -95 156 -89
rect 180 -91 186 -89
rect 137 -103 156 -95
rect 152 -110 156 -103
rect 164 -110 172 -91
rect 180 -103 184 -91
rect 195 -93 201 -91
rect 193 -101 201 -93
rect 195 -103 201 -101
rect 180 -108 186 -103
rect 180 -109 192 -108
rect 180 -110 193 -109
rect 199 -110 201 -108
rect 0 -118 186 -110
rect 190 -111 201 -110
rect 191 -112 201 -111
rect 209 -110 215 -85
rect 223 -110 225 -85
rect 234 -87 238 -85
rect 246 -87 260 -85
rect 270 -87 393 -85
rect 248 -89 258 -87
rect 250 -91 256 -89
rect 264 -91 266 -89
rect 275 -91 393 -87
rect 234 -110 242 -91
rect 250 -103 254 -91
rect 262 -95 268 -91
rect 272 -99 275 -97
rect 277 -99 393 -91
rect 260 -101 393 -99
rect 264 -103 275 -101
rect 250 -106 256 -103
rect 250 -108 258 -106
rect 277 -108 393 -101
rect 250 -110 260 -108
rect 275 -110 393 -108
rect 209 -112 393 -110
rect 207 -114 393 -112
rect 205 -116 393 -114
rect 201 -118 393 -116
rect 0 -124 393 -118
rect 0 -435 35 -124
rect 51 -142 59 -134
rect 98 -136 100 -134
rect 102 -136 104 -134
rect 123 -136 127 -134
rect 133 -136 150 -134
rect 154 -136 156 -134
rect 170 -136 172 -134
rect 64 -138 68 -136
rect 80 -138 84 -136
rect 109 -138 121 -136
rect 133 -138 178 -136
rect 182 -138 184 -136
rect 186 -138 188 -134
rect 193 -136 199 -134
rect 201 -136 205 -134
rect 209 -136 213 -134
rect 217 -136 221 -134
rect 232 -136 238 -134
rect 242 -136 258 -134
rect 262 -136 266 -134
rect 281 -136 285 -134
rect 287 -136 295 -134
rect 299 -136 303 -134
rect 311 -136 315 -134
rect 318 -136 324 -134
rect 191 -138 234 -136
rect 240 -138 248 -136
rect 66 -140 68 -138
rect 74 -140 76 -138
rect 82 -140 84 -138
rect 94 -140 106 -138
rect 109 -140 113 -138
rect 51 -144 53 -142
rect 57 -144 59 -142
rect 64 -144 68 -140
rect 78 -144 80 -142
rect 86 -144 88 -140
rect 94 -142 100 -140
rect 104 -142 113 -140
rect 115 -140 123 -138
rect 133 -140 164 -138
rect 166 -140 238 -138
rect 242 -140 248 -138
rect 252 -138 268 -136
rect 273 -138 277 -136
rect 281 -138 289 -136
rect 291 -138 295 -136
rect 252 -140 266 -138
rect 270 -140 275 -138
rect 281 -140 287 -138
rect 291 -140 297 -138
rect 301 -140 307 -136
rect 309 -138 315 -136
rect 320 -138 326 -136
rect 318 -140 326 -138
rect 328 -140 342 -134
rect 115 -142 119 -140
rect 133 -142 135 -140
rect 139 -142 258 -140
rect 98 -144 100 -142
rect 102 -144 121 -142
rect 139 -144 141 -142
rect 145 -144 168 -142
rect 172 -144 174 -142
rect 178 -144 258 -142
rect 260 -142 266 -140
rect 268 -142 272 -140
rect 279 -142 283 -140
rect 260 -144 264 -142
rect 268 -144 270 -142
rect 275 -144 283 -142
rect 285 -142 295 -140
rect 285 -144 287 -142
rect 293 -144 297 -142
rect 51 -147 66 -144
rect 51 -149 59 -147
rect 64 -149 66 -147
rect 76 -147 82 -144
rect 96 -147 104 -144
rect 107 -147 119 -144
rect 125 -147 129 -144
rect 131 -147 133 -144
rect 76 -149 78 -147
rect 90 -149 94 -147
rect 98 -149 111 -147
rect 113 -149 135 -147
rect 141 -149 145 -147
rect 158 -149 168 -144
rect 184 -147 266 -144
rect 272 -147 277 -144
rect 281 -147 289 -144
rect 295 -147 299 -144
rect 303 -147 307 -140
rect 315 -142 326 -140
rect 332 -142 336 -140
rect 338 -142 342 -140
rect 316 -144 320 -142
rect 324 -144 330 -142
rect 332 -144 342 -142
rect 315 -147 318 -144
rect 322 -147 326 -144
rect 328 -147 342 -144
rect 170 -149 172 -147
rect 191 -149 193 -147
rect 195 -149 205 -147
rect 51 -151 61 -149
rect 86 -151 162 -149
rect 164 -151 178 -149
rect 199 -151 205 -149
rect 207 -149 229 -147
rect 231 -149 252 -147
rect 256 -149 291 -147
rect 313 -149 318 -147
rect 332 -149 342 -147
rect 207 -151 209 -149
rect 223 -151 262 -149
rect 264 -151 272 -149
rect 275 -151 285 -149
rect 287 -151 295 -149
rect 305 -151 307 -149
rect 313 -151 315 -149
rect 324 -151 342 -149
rect 51 -155 57 -151
rect 70 -153 72 -151
rect 84 -153 92 -151
rect 96 -153 182 -151
rect 193 -153 197 -151
rect 199 -153 209 -151
rect 219 -153 293 -151
rect 297 -153 301 -151
rect 305 -153 315 -151
rect 322 -153 342 -151
rect 61 -155 68 -153
rect 90 -155 94 -153
rect 96 -155 203 -153
rect 207 -155 301 -153
rect 51 -157 59 -155
rect 64 -157 70 -155
rect 78 -157 80 -155
rect 92 -157 301 -155
rect 307 -157 309 -153
rect 322 -155 324 -153
rect 330 -155 342 -153
rect 320 -157 324 -155
rect 334 -157 342 -155
rect 51 -159 53 -157
rect 55 -159 61 -157
rect 64 -159 66 -157
rect 88 -159 90 -157
rect 98 -159 295 -157
rect 299 -159 305 -157
rect 320 -159 322 -157
rect 326 -159 330 -157
rect 51 -161 57 -159
rect 64 -161 68 -159
rect 88 -161 92 -159
rect 98 -161 305 -159
rect 311 -161 313 -159
rect 324 -161 330 -159
rect 332 -159 342 -157
rect 332 -161 338 -159
rect 51 -165 55 -161
rect 59 -163 66 -161
rect 76 -163 82 -161
rect 88 -163 94 -161
rect 102 -163 143 -161
rect 158 -163 299 -161
rect 57 -165 64 -163
rect 80 -165 84 -163
rect 90 -165 94 -163
rect 98 -165 139 -163
rect 53 -167 59 -165
rect 62 -167 66 -165
rect 72 -167 76 -165
rect 92 -167 96 -165
rect 100 -167 107 -165
rect 109 -167 127 -165
rect 129 -167 139 -165
rect 141 -167 143 -163
rect 51 -171 64 -167
rect 74 -169 78 -167
rect 100 -169 125 -167
rect 70 -171 80 -169
rect 100 -171 104 -169
rect 107 -171 125 -169
rect 51 -173 59 -171
rect 61 -173 66 -171
rect 72 -173 74 -171
rect 88 -173 96 -171
rect 51 -175 53 -173
rect 61 -175 68 -173
rect 94 -175 98 -173
rect 102 -175 109 -171
rect 111 -173 125 -171
rect 131 -171 139 -167
rect 148 -169 156 -163
rect 164 -165 299 -163
rect 309 -163 313 -161
rect 332 -163 342 -161
rect 309 -165 311 -163
rect 315 -165 320 -163
rect 330 -165 342 -163
rect 164 -167 246 -165
rect 252 -167 303 -165
rect 313 -167 320 -165
rect 324 -167 328 -165
rect 164 -169 231 -167
rect 141 -171 145 -169
rect 131 -173 145 -171
rect 162 -171 176 -169
rect 180 -171 231 -169
rect 162 -173 178 -171
rect 182 -173 231 -171
rect 234 -169 248 -167
rect 252 -169 254 -167
rect 234 -171 246 -169
rect 250 -171 254 -169
rect 256 -171 297 -167
rect 326 -169 328 -167
rect 332 -169 336 -165
rect 340 -167 342 -165
rect 324 -171 334 -169
rect 338 -171 342 -167
rect 234 -173 238 -171
rect 252 -173 264 -171
rect 268 -173 301 -171
rect 322 -173 328 -171
rect 330 -173 334 -171
rect 336 -173 342 -171
rect 113 -175 125 -173
rect 133 -175 148 -173
rect 156 -175 180 -173
rect 182 -175 236 -173
rect 250 -175 264 -173
rect 51 -177 55 -175
rect 59 -177 64 -175
rect 66 -177 72 -175
rect 86 -177 88 -175
rect 107 -177 111 -175
rect 113 -177 129 -175
rect 51 -179 68 -177
rect 70 -179 72 -177
rect 107 -179 129 -177
rect 135 -179 172 -175
rect 174 -177 180 -175
rect 184 -177 238 -175
rect 246 -177 264 -175
rect 174 -179 264 -177
rect 270 -175 287 -173
rect 291 -175 293 -173
rect 295 -175 299 -173
rect 270 -179 283 -175
rect 291 -177 297 -175
rect 318 -177 324 -173
rect 330 -175 340 -173
rect 328 -177 340 -175
rect 289 -179 293 -177
rect 303 -179 307 -177
rect 328 -179 342 -177
rect 51 -181 57 -179
rect 64 -181 66 -179
rect 104 -181 131 -179
rect 135 -181 137 -179
rect 141 -181 213 -179
rect 219 -181 262 -179
rect 270 -181 281 -179
rect 285 -181 293 -179
rect 297 -181 301 -179
rect 303 -181 305 -179
rect 326 -181 330 -179
rect 332 -181 334 -179
rect 338 -181 342 -179
rect 51 -183 55 -181
rect 59 -183 61 -181
rect 78 -183 80 -181
rect 104 -183 109 -181
rect 111 -183 133 -181
rect 145 -183 168 -181
rect 170 -183 174 -181
rect 176 -183 217 -181
rect 227 -183 260 -181
rect 264 -183 281 -181
rect 287 -183 291 -181
rect 51 -185 53 -183
rect 57 -185 61 -183
rect 96 -185 98 -183
rect 107 -185 135 -183
rect 148 -185 166 -183
rect 172 -185 221 -183
rect 229 -185 260 -183
rect 262 -185 281 -183
rect 51 -190 55 -185
rect 57 -187 59 -185
rect 100 -187 102 -185
rect 107 -187 139 -185
rect 154 -187 158 -185
rect 160 -187 166 -185
rect 168 -187 281 -185
rect 283 -185 293 -183
rect 303 -185 307 -183
rect 315 -185 320 -181
rect 326 -183 334 -181
rect 283 -187 285 -185
rect 289 -187 295 -185
rect 303 -187 305 -185
rect 57 -190 61 -187
rect 90 -190 92 -187
rect 104 -190 113 -187
rect 117 -190 121 -187
rect 123 -190 145 -187
rect 154 -190 184 -187
rect 186 -190 229 -187
rect 234 -190 238 -187
rect 242 -190 246 -187
rect 51 -194 53 -190
rect 76 -194 78 -190
rect 94 -192 98 -190
rect 104 -192 115 -190
rect 117 -192 182 -190
rect 186 -192 197 -190
rect 94 -194 96 -192
rect 111 -194 154 -192
rect 170 -194 182 -192
rect 51 -198 55 -194
rect 59 -196 66 -194
rect 109 -196 115 -194
rect 119 -196 145 -194
rect 174 -196 182 -194
rect 184 -194 197 -192
rect 184 -196 188 -194
rect 191 -196 197 -194
rect 57 -198 61 -196
rect 109 -198 131 -196
rect 133 -198 145 -196
rect 176 -198 197 -196
rect 51 -200 66 -198
rect 109 -200 111 -198
rect 113 -200 154 -198
rect 174 -200 186 -198
rect 51 -202 53 -200
rect 55 -202 57 -200
rect 61 -202 66 -200
rect 94 -202 98 -200
rect 104 -202 107 -200
rect 113 -202 143 -200
rect 176 -202 186 -200
rect 188 -202 197 -198
rect 51 -206 59 -202
rect 64 -204 74 -202
rect 102 -204 109 -202
rect 111 -204 115 -202
rect 117 -204 141 -202
rect 68 -206 70 -204
rect 94 -206 96 -204
rect 102 -206 104 -204
rect 107 -206 143 -204
rect 176 -206 184 -202
rect 188 -204 193 -202
rect 195 -204 197 -202
rect 199 -192 236 -190
rect 240 -192 246 -190
rect 250 -190 277 -187
rect 279 -190 291 -187
rect 324 -190 328 -183
rect 336 -187 342 -181
rect 332 -190 338 -187
rect 250 -192 264 -190
rect 268 -192 283 -190
rect 285 -192 291 -190
rect 199 -194 264 -192
rect 266 -194 281 -192
rect 297 -194 303 -190
rect 309 -192 311 -190
rect 324 -192 330 -190
rect 334 -192 342 -190
rect 309 -194 315 -192
rect 326 -194 332 -192
rect 199 -196 281 -194
rect 283 -196 287 -194
rect 328 -196 332 -194
rect 199 -198 209 -196
rect 213 -198 223 -196
rect 231 -198 289 -196
rect 199 -200 207 -198
rect 211 -200 221 -198
rect 246 -200 283 -198
rect 293 -200 299 -198
rect 305 -200 309 -196
rect 315 -198 324 -196
rect 328 -198 330 -196
rect 336 -198 342 -192
rect 315 -200 320 -198
rect 326 -200 342 -198
rect 199 -204 209 -200
rect 186 -206 193 -204
rect 55 -208 59 -206
rect 94 -208 98 -206
rect 102 -208 145 -206
rect 55 -210 61 -208
rect 107 -210 109 -208
rect 111 -210 133 -208
rect 148 -210 150 -208
rect 51 -214 57 -210
rect 59 -212 61 -210
rect 66 -212 70 -210
rect 100 -212 104 -210
rect 107 -212 133 -210
rect 98 -214 102 -212
rect 109 -214 113 -212
rect 115 -214 123 -212
rect 125 -214 133 -212
rect 51 -216 55 -214
rect 61 -216 66 -214
rect 90 -216 92 -214
rect 104 -216 121 -214
rect 125 -216 139 -214
rect 51 -220 57 -216
rect 64 -220 68 -216
rect 102 -218 107 -216
rect 109 -218 117 -216
rect 119 -218 133 -216
rect 137 -218 141 -216
rect 178 -218 182 -206
rect 186 -208 195 -206
rect 201 -208 209 -204
rect 213 -204 219 -200
rect 248 -202 283 -200
rect 297 -202 301 -200
rect 307 -202 309 -200
rect 313 -202 318 -200
rect 328 -202 336 -200
rect 340 -202 342 -200
rect 244 -204 281 -202
rect 186 -212 193 -208
rect 201 -210 207 -208
rect 199 -212 209 -210
rect 213 -212 221 -204
rect 242 -206 248 -204
rect 252 -206 281 -204
rect 287 -206 295 -202
rect 326 -204 336 -202
rect 301 -206 305 -204
rect 318 -206 320 -204
rect 324 -206 328 -204
rect 330 -206 342 -204
rect 240 -208 244 -206
rect 254 -210 277 -206
rect 279 -208 285 -206
rect 291 -208 293 -206
rect 301 -208 313 -206
rect 318 -208 342 -206
rect 281 -210 289 -208
rect 291 -210 295 -208
rect 303 -210 305 -208
rect 311 -210 313 -208
rect 320 -210 324 -208
rect 254 -212 287 -210
rect 199 -214 211 -212
rect 186 -216 188 -214
rect 191 -218 193 -216
rect 199 -218 209 -214
rect 102 -220 104 -218
rect 115 -220 117 -218
rect 121 -220 131 -218
rect 139 -220 143 -218
rect 51 -222 55 -220
rect 64 -222 70 -220
rect 113 -222 131 -220
rect 141 -222 143 -220
rect 51 -224 57 -222
rect 104 -224 109 -222
rect 113 -224 115 -222
rect 117 -224 121 -222
rect 123 -224 129 -222
rect 51 -226 66 -224
rect 104 -226 107 -224
rect 55 -228 66 -226
rect 86 -228 88 -226
rect 119 -228 121 -226
rect 125 -228 129 -224
rect 178 -226 180 -218
rect 191 -220 195 -218
rect 201 -222 211 -218
rect 215 -220 221 -212
rect 252 -214 256 -212
rect 260 -214 287 -212
rect 293 -212 299 -210
rect 307 -212 318 -210
rect 322 -212 324 -210
rect 326 -210 330 -208
rect 332 -210 342 -208
rect 326 -212 342 -210
rect 293 -214 301 -212
rect 305 -214 311 -212
rect 315 -214 320 -212
rect 322 -214 330 -212
rect 334 -214 342 -212
rect 197 -224 199 -222
rect 203 -226 211 -222
rect 217 -226 221 -220
rect 51 -231 57 -228
rect 64 -230 68 -228
rect 117 -230 121 -228
rect 123 -230 129 -228
rect 51 -233 59 -231
rect 117 -233 129 -230
rect 51 -235 55 -233
rect 57 -235 61 -233
rect 113 -235 127 -233
rect 178 -235 180 -228
rect 186 -235 188 -230
rect 195 -233 197 -228
rect 205 -230 211 -226
rect 207 -235 211 -230
rect 51 -239 64 -235
rect 68 -237 72 -235
rect 111 -237 117 -235
rect 119 -237 125 -235
rect 68 -239 82 -237
rect 111 -239 125 -237
rect 51 -241 66 -239
rect 68 -241 72 -239
rect 102 -241 104 -239
rect 109 -241 113 -239
rect 51 -243 59 -241
rect 64 -243 72 -241
rect 100 -243 104 -241
rect 107 -243 111 -241
rect 119 -243 125 -239
rect 178 -237 182 -235
rect 51 -247 66 -243
rect 68 -245 74 -243
rect 102 -245 109 -243
rect 121 -245 123 -243
rect 70 -247 72 -245
rect 51 -249 72 -247
rect 51 -251 64 -249
rect 68 -251 72 -249
rect 78 -247 84 -245
rect 90 -247 92 -245
rect 104 -247 109 -245
rect 117 -247 125 -245
rect 78 -249 80 -247
rect 82 -249 84 -247
rect 107 -249 113 -247
rect 78 -251 84 -249
rect 109 -251 113 -249
rect 115 -251 125 -247
rect 178 -249 180 -237
rect 186 -239 188 -237
rect 205 -239 211 -235
rect 219 -237 221 -226
rect 262 -218 275 -214
rect 277 -216 289 -214
rect 295 -216 297 -214
rect 305 -216 313 -214
rect 324 -216 342 -214
rect 279 -218 293 -216
rect 295 -218 299 -216
rect 305 -218 309 -216
rect 311 -218 313 -216
rect 318 -218 322 -216
rect 324 -218 338 -216
rect 262 -220 277 -218
rect 285 -220 299 -218
rect 307 -220 342 -218
rect 262 -224 283 -220
rect 303 -222 305 -220
rect 307 -222 316 -220
rect 320 -222 326 -220
rect 289 -224 293 -222
rect 295 -224 299 -222
rect 309 -224 313 -222
rect 318 -224 322 -222
rect 328 -224 342 -220
rect 262 -226 272 -224
rect 275 -226 285 -224
rect 289 -226 299 -224
rect 305 -226 311 -224
rect 315 -226 320 -224
rect 324 -226 334 -224
rect 336 -226 342 -224
rect 262 -228 277 -226
rect 266 -230 277 -228
rect 279 -228 287 -226
rect 301 -228 309 -226
rect 279 -230 293 -228
rect 266 -233 285 -230
rect 287 -233 293 -230
rect 299 -230 309 -228
rect 313 -228 342 -226
rect 313 -230 322 -228
rect 324 -230 342 -228
rect 299 -233 305 -230
rect 307 -233 328 -230
rect 330 -233 342 -230
rect 260 -235 262 -233
rect 266 -235 279 -233
rect 281 -235 285 -233
rect 299 -235 313 -233
rect 315 -235 342 -233
rect 266 -239 285 -235
rect 287 -237 289 -235
rect 303 -237 305 -235
rect 309 -237 313 -235
rect 320 -237 342 -235
rect 303 -239 315 -237
rect 324 -239 342 -237
rect 205 -245 213 -239
rect 219 -243 221 -239
rect 268 -241 291 -239
rect 297 -241 299 -239
rect 307 -241 309 -239
rect 313 -241 320 -239
rect 268 -243 293 -241
rect 295 -243 301 -241
rect 311 -243 324 -241
rect 326 -243 342 -239
rect 184 -247 190 -245
rect 188 -249 191 -247
rect 207 -249 213 -245
rect 268 -247 281 -243
rect 285 -245 299 -243
rect 307 -245 342 -243
rect 283 -247 293 -245
rect 305 -247 342 -245
rect 268 -249 279 -247
rect 285 -249 287 -247
rect 178 -251 182 -249
rect 207 -251 215 -249
rect 270 -251 281 -249
rect 291 -251 295 -249
rect 301 -251 307 -247
rect 309 -249 332 -247
rect 313 -251 332 -249
rect 334 -251 342 -247
rect 51 -253 74 -251
rect 76 -253 88 -251
rect 92 -253 94 -251
rect 100 -253 104 -251
rect 111 -253 125 -251
rect 209 -253 213 -251
rect 270 -253 289 -251
rect 293 -253 295 -251
rect 303 -253 311 -251
rect 51 -255 72 -253
rect 78 -255 84 -253
rect 98 -255 104 -253
rect 109 -255 125 -253
rect 51 -257 55 -255
rect 57 -257 76 -255
rect 82 -257 86 -255
rect 51 -259 68 -257
rect 72 -259 78 -257
rect 84 -259 90 -257
rect 98 -259 100 -257
rect 51 -263 78 -259
rect 80 -263 84 -261
rect 86 -263 88 -259
rect 94 -261 96 -259
rect 104 -261 109 -259
rect 111 -261 127 -255
rect 207 -257 213 -253
rect 272 -255 285 -253
rect 287 -255 291 -253
rect 297 -255 305 -253
rect 307 -255 311 -253
rect 313 -255 342 -251
rect 272 -257 291 -255
rect 299 -257 342 -255
rect 178 -259 182 -257
rect 184 -259 186 -257
rect 188 -259 191 -257
rect 207 -259 215 -257
rect 104 -263 127 -261
rect 51 -265 92 -263
rect 96 -265 100 -263
rect 104 -265 111 -263
rect 113 -265 127 -263
rect 180 -261 182 -259
rect 188 -261 193 -259
rect 205 -261 215 -259
rect 272 -261 289 -257
rect 293 -259 301 -257
rect 305 -259 334 -257
rect 336 -259 342 -257
rect 291 -261 303 -259
rect 305 -261 340 -259
rect 180 -265 184 -261
rect 188 -263 191 -261
rect 205 -263 213 -261
rect 51 -269 53 -265
rect 57 -267 70 -265
rect 74 -267 82 -265
rect 86 -267 92 -265
rect 94 -267 107 -265
rect 55 -269 90 -267
rect 98 -269 104 -267
rect 109 -269 111 -267
rect 113 -269 129 -265
rect 51 -271 94 -269
rect 96 -271 129 -269
rect 51 -274 84 -271
rect 88 -272 98 -271
rect 90 -274 98 -272
rect 51 -276 88 -274
rect 92 -276 96 -274
rect 100 -276 129 -271
rect 51 -284 129 -276
rect 180 -267 182 -265
rect 207 -267 211 -263
rect 264 -265 266 -261
rect 213 -267 215 -265
rect 180 -271 186 -267
rect 205 -269 215 -267
rect 221 -269 223 -265
rect 262 -267 266 -265
rect 270 -263 340 -261
rect 270 -265 332 -263
rect 334 -265 342 -263
rect 205 -271 217 -269
rect 180 -274 184 -271
rect 205 -274 207 -271
rect 215 -274 217 -271
rect 262 -272 264 -267
rect 260 -274 264 -272
rect 270 -269 297 -265
rect 299 -269 342 -265
rect 270 -271 340 -269
rect 270 -274 342 -271
rect 180 -278 186 -274
rect 195 -278 197 -276
rect 205 -278 213 -274
rect 180 -282 184 -278
rect 182 -284 184 -282
rect 188 -280 193 -278
rect 188 -284 191 -280
rect 205 -282 215 -278
rect 219 -280 223 -274
rect 260 -278 262 -274
rect 270 -278 332 -274
rect 338 -276 342 -274
rect 336 -278 342 -276
rect 268 -280 330 -278
rect 334 -280 340 -278
rect 221 -282 223 -280
rect 209 -284 215 -282
rect 51 -286 88 -284
rect 90 -286 107 -284
rect 109 -286 131 -284
rect 51 -288 113 -286
rect 115 -288 131 -286
rect 182 -286 193 -284
rect 209 -286 217 -284
rect 219 -286 221 -284
rect 258 -286 260 -280
rect 268 -282 322 -280
rect 324 -282 328 -280
rect 268 -284 320 -282
rect 324 -284 326 -282
rect 334 -284 336 -280
rect 182 -288 188 -286
rect 207 -288 221 -286
rect 266 -288 320 -284
rect 322 -286 326 -284
rect 324 -288 326 -286
rect 51 -296 133 -288
rect 182 -292 184 -288
rect 186 -290 193 -288
rect 188 -292 193 -290
rect 203 -290 205 -288
rect 207 -290 219 -288
rect 203 -292 213 -290
rect 256 -292 258 -288
rect 266 -292 307 -288
rect 182 -294 191 -292
rect 205 -294 215 -292
rect 264 -294 311 -292
rect 51 -298 135 -296
rect 51 -300 90 -298
rect 92 -300 135 -298
rect 51 -302 135 -300
rect 184 -300 193 -294
rect 201 -296 213 -294
rect 264 -296 318 -294
rect 203 -298 219 -296
rect 262 -298 322 -296
rect 184 -302 197 -300
rect 199 -302 201 -300
rect 205 -302 217 -298
rect 262 -300 320 -298
rect 252 -302 254 -300
rect 262 -302 315 -300
rect 51 -306 137 -302
rect 186 -304 197 -302
rect 143 -306 145 -304
rect 51 -308 86 -306
rect 88 -308 137 -306
rect 160 -308 162 -304
rect 51 -310 139 -308
rect 145 -310 148 -308
rect 160 -310 164 -308
rect 174 -310 176 -306
rect 186 -308 193 -304
rect 203 -308 217 -302
rect 260 -304 315 -302
rect 322 -304 324 -300
rect 260 -306 309 -304
rect 313 -306 318 -304
rect 258 -308 322 -306
rect 186 -310 191 -308
rect 203 -310 219 -308
rect 51 -312 141 -310
rect 145 -312 150 -310
rect 51 -314 96 -312
rect 98 -314 137 -312
rect 51 -315 137 -314
rect 139 -314 141 -312
rect 148 -314 152 -312
rect 139 -315 143 -314
rect 51 -317 143 -315
rect 150 -317 152 -314
rect 162 -314 164 -310
rect 51 -319 139 -317
rect 141 -319 145 -317
rect 150 -319 154 -317
rect 162 -319 166 -314
rect 51 -321 145 -319
rect 152 -321 154 -319
rect 158 -321 160 -319
rect 162 -321 168 -319
rect 51 -323 133 -321
rect 135 -323 141 -321
rect 143 -323 148 -321
rect 152 -323 156 -321
rect 164 -323 168 -321
rect 176 -321 178 -312
rect 186 -317 188 -310
rect 207 -312 219 -310
rect 238 -312 240 -310
rect 258 -312 260 -308
rect 262 -312 318 -308
rect 195 -314 197 -312
rect 203 -314 205 -312
rect 207 -317 217 -312
rect 236 -314 240 -312
rect 248 -314 250 -312
rect 256 -314 324 -312
rect 221 -317 223 -314
rect 236 -317 238 -314
rect 246 -317 250 -314
rect 254 -317 309 -314
rect 315 -317 324 -314
rect 184 -319 190 -317
rect 207 -319 219 -317
rect 176 -323 180 -321
rect 184 -323 186 -319
rect 188 -321 191 -319
rect 207 -321 221 -319
rect 236 -321 240 -317
rect 244 -319 248 -317
rect 254 -319 256 -317
rect 258 -319 309 -317
rect 322 -319 326 -317
rect 195 -323 199 -321
rect 207 -323 223 -321
rect 51 -325 141 -323
rect 145 -325 150 -323
rect 51 -329 143 -325
rect 145 -327 152 -325
rect 154 -327 156 -323
rect 166 -325 168 -323
rect 178 -325 182 -323
rect 207 -325 219 -323
rect 148 -329 164 -327
rect 51 -331 145 -329
rect 51 -333 148 -331
rect 150 -333 154 -329
rect 156 -333 160 -329
rect 162 -331 164 -329
rect 166 -331 170 -325
rect 191 -327 195 -325
rect 199 -327 201 -325
rect 209 -327 211 -325
rect 215 -327 219 -325
rect 221 -327 223 -323
rect 182 -329 184 -327
rect 193 -329 195 -327
rect 215 -329 223 -327
rect 234 -327 238 -321
rect 242 -323 248 -319
rect 252 -321 318 -319
rect 324 -321 328 -319
rect 252 -323 311 -321
rect 315 -323 318 -321
rect 326 -323 328 -321
rect 244 -325 248 -323
rect 250 -325 254 -323
rect 258 -325 311 -323
rect 244 -327 252 -325
rect 234 -329 252 -327
rect 256 -327 277 -325
rect 256 -329 281 -327
rect 283 -329 311 -325
rect 209 -331 221 -329
rect 242 -331 311 -329
rect 178 -333 180 -331
rect 211 -333 215 -331
rect 217 -333 225 -331
rect 227 -333 233 -331
rect 244 -333 277 -331
rect 289 -333 295 -331
rect 297 -333 315 -331
rect 51 -335 125 -333
rect 127 -335 154 -333
rect 158 -335 160 -333
rect 174 -335 186 -333
rect 219 -335 225 -333
rect 231 -335 236 -333
rect 240 -335 277 -333
rect 293 -335 311 -333
rect 51 -337 115 -335
rect 117 -337 150 -335
rect 152 -337 160 -335
rect 170 -337 172 -335
rect 191 -337 193 -335
rect 217 -337 221 -335
rect 231 -337 234 -335
rect 51 -339 156 -337
rect 158 -339 166 -337
rect 191 -339 195 -337
rect 219 -339 225 -337
rect 242 -339 275 -335
rect 295 -337 311 -335
rect 313 -337 315 -333
rect 295 -339 315 -337
rect 51 -341 98 -339
rect 100 -341 154 -339
rect 160 -341 164 -339
rect 201 -341 203 -339
rect 223 -341 225 -339
rect 240 -341 244 -339
rect 248 -341 275 -339
rect 51 -343 86 -341
rect 92 -343 162 -341
rect 186 -343 191 -341
rect 215 -343 219 -341
rect 238 -343 244 -341
rect 246 -343 272 -341
rect 51 -345 84 -343
rect 88 -345 111 -343
rect 117 -345 133 -343
rect 51 -347 57 -345
rect 59 -347 133 -345
rect 135 -347 143 -343
rect 51 -349 123 -347
rect 127 -349 143 -347
rect 145 -347 152 -343
rect 154 -345 160 -343
rect 231 -345 248 -343
rect 250 -345 270 -343
rect 154 -347 158 -345
rect 145 -349 158 -347
rect 172 -347 180 -345
rect 227 -347 246 -345
rect 250 -347 272 -345
rect 297 -347 313 -339
rect 172 -349 186 -347
rect 225 -349 238 -347
rect 248 -349 272 -347
rect 51 -351 55 -349
rect 57 -351 102 -349
rect 107 -351 111 -349
rect 115 -351 117 -349
rect 119 -351 123 -349
rect 125 -351 143 -349
rect 148 -351 158 -349
rect 170 -351 188 -349
rect 223 -351 234 -349
rect 242 -351 272 -349
rect 295 -349 311 -347
rect 295 -351 301 -349
rect 51 -358 53 -351
rect 59 -353 96 -351
rect 115 -353 143 -351
rect 145 -353 156 -351
rect 180 -353 191 -351
rect 221 -353 229 -351
rect 240 -353 244 -351
rect 248 -353 268 -351
rect 297 -353 301 -351
rect 303 -351 311 -349
rect 303 -353 313 -351
rect 57 -355 68 -353
rect 70 -355 94 -353
rect 104 -355 107 -353
rect 113 -355 125 -353
rect 127 -355 139 -353
rect 141 -355 158 -353
rect 186 -355 193 -353
rect 219 -355 227 -353
rect 234 -355 238 -353
rect 242 -355 270 -353
rect 57 -358 88 -355
rect 111 -358 117 -355
rect 119 -358 145 -355
rect 148 -358 158 -355
rect 188 -358 195 -355
rect 219 -358 225 -355
rect 244 -358 272 -355
rect 293 -358 295 -353
rect 299 -355 309 -353
rect 299 -358 311 -355
rect 55 -360 86 -358
rect 119 -360 158 -358
rect 191 -360 195 -358
rect 217 -360 223 -358
rect 242 -360 268 -358
rect 301 -360 309 -358
rect 55 -362 78 -360
rect 80 -362 94 -360
rect 115 -362 158 -360
rect 178 -362 180 -360
rect 193 -362 197 -360
rect 215 -362 221 -360
rect 248 -362 264 -360
rect 266 -362 270 -360
rect 59 -364 88 -362
rect 111 -364 117 -362
rect 119 -364 135 -362
rect 137 -364 158 -362
rect 195 -364 199 -362
rect 57 -366 61 -364
rect 70 -366 84 -364
rect 111 -366 113 -364
rect 123 -366 129 -364
rect 133 -366 158 -364
rect 160 -366 162 -364
rect 197 -366 201 -364
rect 213 -366 219 -362
rect 248 -364 260 -362
rect 289 -364 291 -360
rect 295 -364 299 -360
rect 301 -362 311 -360
rect 303 -364 311 -362
rect 221 -366 223 -364
rect 246 -366 262 -364
rect 297 -366 301 -364
rect 57 -368 59 -366
rect 66 -368 84 -366
rect 115 -368 117 -366
rect 123 -368 127 -366
rect 133 -368 162 -366
rect 199 -368 201 -366
rect 227 -368 229 -366
rect 231 -368 238 -366
rect 240 -368 242 -366
rect 64 -370 86 -368
rect 113 -370 119 -368
rect 131 -370 158 -368
rect 160 -370 164 -368
rect 213 -370 215 -368
rect 231 -370 242 -368
rect 246 -368 264 -366
rect 287 -368 289 -366
rect 291 -368 295 -366
rect 246 -370 254 -368
rect 268 -370 270 -368
rect 293 -370 295 -368
rect 299 -370 301 -366
rect 303 -366 309 -364
rect 303 -368 307 -366
rect 61 -372 88 -370
rect 64 -374 88 -372
rect 117 -374 123 -370
rect 131 -372 137 -370
rect 141 -372 150 -370
rect 154 -372 166 -370
rect 186 -372 188 -370
rect 197 -372 199 -370
rect 131 -374 135 -372
rect 139 -374 148 -372
rect 152 -374 164 -372
rect 203 -374 205 -370
rect 213 -372 217 -370
rect 225 -372 229 -370
rect 231 -372 240 -370
rect 244 -372 258 -370
rect 268 -372 272 -370
rect 275 -372 281 -370
rect 297 -372 303 -370
rect 305 -372 309 -368
rect 213 -374 215 -372
rect 223 -374 227 -372
rect 234 -374 236 -372
rect 242 -374 254 -372
rect 256 -374 258 -372
rect 270 -374 272 -372
rect 279 -374 283 -372
rect 295 -374 299 -372
rect 57 -376 59 -374
rect 55 -378 61 -376
rect 64 -378 86 -374
rect 115 -376 121 -374
rect 131 -376 133 -374
rect 137 -376 148 -374
rect 150 -376 154 -374
rect 115 -378 119 -376
rect 129 -378 133 -376
rect 139 -378 145 -376
rect 150 -378 152 -376
rect 156 -378 160 -374
rect 166 -376 168 -374
rect 203 -376 207 -374
rect 211 -376 215 -374
rect 162 -378 168 -376
rect 170 -378 172 -376
rect 205 -378 207 -376
rect 209 -378 215 -376
rect 225 -376 227 -374
rect 231 -376 240 -374
rect 248 -376 254 -374
rect 225 -378 242 -376
rect 250 -378 252 -376
rect 266 -378 268 -374
rect 281 -376 285 -374
rect 291 -376 293 -374
rect 283 -378 285 -376
rect 55 -382 57 -378
rect 64 -380 84 -378
rect 127 -380 133 -378
rect 148 -380 152 -378
rect 154 -380 174 -378
rect 197 -380 201 -378
rect 68 -382 84 -380
rect 125 -382 131 -380
rect 137 -382 139 -380
rect 148 -382 150 -380
rect 158 -382 170 -380
rect 172 -382 174 -380
rect 178 -382 182 -380
rect 184 -382 186 -380
rect 59 -384 64 -382
rect 68 -384 80 -382
rect 123 -384 129 -382
rect 133 -384 139 -382
rect 156 -384 162 -382
rect 166 -384 168 -382
rect 172 -384 176 -382
rect 180 -384 182 -382
rect 199 -384 201 -380
rect 205 -380 215 -378
rect 223 -380 227 -378
rect 231 -380 234 -378
rect 236 -380 244 -378
rect 287 -380 293 -376
rect 297 -380 299 -374
rect 301 -376 303 -372
rect 307 -376 309 -372
rect 205 -382 219 -380
rect 223 -382 229 -380
rect 231 -382 238 -380
rect 242 -382 246 -380
rect 260 -382 262 -380
rect 285 -382 293 -380
rect 51 -386 53 -384
rect 57 -386 64 -384
rect 66 -386 80 -384
rect 86 -386 92 -384
rect 123 -386 137 -384
rect 156 -386 160 -384
rect 164 -386 168 -384
rect 170 -386 174 -384
rect 184 -386 186 -384
rect 51 -388 55 -386
rect 57 -388 61 -386
rect 51 -390 61 -388
rect 66 -388 92 -386
rect 96 -388 104 -386
rect 119 -388 121 -386
rect 66 -390 90 -388
rect 117 -390 121 -388
rect 129 -388 137 -386
rect 164 -388 166 -386
rect 170 -388 172 -386
rect 176 -388 180 -386
rect 182 -388 188 -386
rect 51 -392 59 -390
rect 64 -392 88 -390
rect 55 -394 57 -392
rect 53 -396 57 -394
rect 61 -394 88 -392
rect 92 -394 94 -390
rect 129 -392 135 -388
rect 139 -390 141 -388
rect 145 -392 148 -388
rect 168 -390 172 -388
rect 174 -390 188 -388
rect 191 -390 195 -384
rect 197 -390 201 -384
rect 203 -384 215 -382
rect 203 -386 205 -384
rect 209 -386 215 -384
rect 217 -384 221 -382
rect 223 -384 236 -382
rect 258 -384 264 -382
rect 285 -384 295 -382
rect 299 -384 301 -382
rect 217 -386 231 -384
rect 234 -386 236 -384
rect 238 -386 240 -384
rect 260 -386 262 -384
rect 270 -386 272 -384
rect 203 -388 207 -386
rect 213 -388 225 -386
rect 203 -390 209 -388
rect 213 -390 215 -388
rect 227 -390 231 -386
rect 287 -388 295 -384
rect 297 -386 301 -384
rect 297 -388 299 -386
rect 307 -388 309 -386
rect 256 -390 260 -388
rect 285 -390 289 -388
rect 297 -390 301 -388
rect 168 -392 170 -390
rect 174 -392 178 -390
rect 182 -392 186 -390
rect 191 -392 193 -390
rect 203 -392 205 -390
rect 258 -392 262 -390
rect 285 -392 291 -390
rect 293 -392 295 -390
rect 299 -392 303 -390
rect 305 -392 309 -390
rect 61 -396 64 -394
rect 66 -396 94 -394
rect 98 -396 100 -394
rect 115 -396 117 -392
rect 125 -394 131 -392
rect 133 -394 137 -392
rect 143 -394 148 -392
rect 184 -394 186 -392
rect 277 -394 281 -392
rect 289 -394 291 -392
rect 125 -396 129 -394
rect 135 -396 137 -394
rect 141 -396 145 -394
rect 244 -396 248 -394
rect 279 -396 281 -394
rect 283 -396 285 -394
rect 289 -396 293 -394
rect 301 -396 303 -392
rect 307 -394 309 -392
rect 51 -398 57 -396
rect 59 -398 100 -396
rect 102 -398 107 -396
rect 125 -398 127 -396
rect 131 -398 137 -396
rect 51 -401 55 -398
rect 59 -401 96 -398
rect 129 -401 135 -398
rect 139 -399 145 -396
rect 152 -398 154 -396
rect 244 -398 250 -396
rect 270 -398 272 -396
rect 279 -398 287 -396
rect 139 -401 147 -399
rect 150 -401 154 -398
rect 158 -401 160 -398
rect 51 -403 57 -401
rect 59 -403 98 -401
rect 51 -405 98 -403
rect 100 -405 104 -403
rect 125 -405 127 -403
rect 131 -405 133 -401
rect 137 -403 143 -401
rect 145 -403 160 -401
rect 164 -403 166 -398
rect 172 -399 174 -398
rect 170 -401 174 -399
rect 207 -401 209 -398
rect 217 -401 219 -398
rect 227 -401 229 -398
rect 275 -401 277 -398
rect 283 -401 287 -398
rect 170 -403 172 -401
rect 205 -403 209 -401
rect 211 -403 213 -401
rect 215 -403 219 -401
rect 223 -403 225 -401
rect 137 -405 141 -403
rect 148 -405 150 -403
rect 154 -405 158 -403
rect 51 -407 111 -405
rect 51 -411 68 -407
rect 70 -411 111 -407
rect 135 -409 141 -405
rect 145 -409 150 -405
rect 152 -407 158 -405
rect 162 -405 166 -403
rect 162 -407 164 -405
rect 168 -407 172 -403
rect 176 -407 178 -403
rect 188 -407 193 -403
rect 201 -407 203 -403
rect 211 -405 227 -403
rect 234 -405 236 -403
rect 268 -405 272 -401
rect 275 -403 279 -401
rect 283 -403 289 -401
rect 291 -403 295 -396
rect 311 -401 313 -398
rect 277 -405 281 -403
rect 285 -405 295 -403
rect 209 -407 219 -405
rect 152 -409 154 -407
rect 166 -409 172 -407
rect 174 -409 178 -407
rect 117 -411 119 -409
rect 51 -413 111 -411
rect 113 -413 119 -411
rect 51 -415 72 -413
rect 76 -415 119 -413
rect 123 -411 127 -409
rect 137 -411 139 -409
rect 145 -411 154 -409
rect 156 -411 160 -409
rect 166 -411 170 -409
rect 174 -411 180 -409
rect 191 -411 197 -407
rect 201 -409 207 -407
rect 209 -409 221 -407
rect 223 -409 227 -405
rect 270 -407 275 -405
rect 279 -407 283 -405
rect 285 -407 291 -405
rect 201 -411 225 -409
rect 270 -411 293 -407
rect 297 -411 301 -409
rect 123 -415 125 -411
rect 148 -413 150 -411
rect 152 -415 158 -411
rect 162 -413 170 -411
rect 172 -413 180 -411
rect 162 -415 164 -413
rect 166 -415 168 -413
rect 172 -415 174 -413
rect 176 -415 180 -413
rect 184 -413 186 -411
rect 191 -413 199 -411
rect 201 -413 223 -411
rect 184 -415 188 -413
rect 191 -415 195 -413
rect 197 -415 199 -413
rect 203 -415 205 -413
rect 207 -415 211 -413
rect 213 -415 219 -413
rect 266 -415 285 -411
rect 287 -415 293 -411
rect 51 -419 74 -415
rect 76 -417 109 -415
rect 111 -417 119 -415
rect 152 -417 156 -415
rect 160 -417 164 -415
rect 178 -417 180 -415
rect 186 -417 188 -415
rect 76 -419 119 -417
rect 51 -421 119 -419
rect 121 -421 123 -417
rect 197 -419 201 -415
rect 266 -417 293 -415
rect 295 -415 297 -413
rect 295 -417 299 -415
rect 334 -417 338 -415
rect 264 -419 289 -417
rect 291 -419 293 -417
rect 258 -421 262 -419
rect 264 -421 293 -419
rect 297 -419 301 -417
rect 311 -419 313 -417
rect 297 -421 303 -419
rect 51 -425 74 -421
rect 76 -425 127 -421
rect 260 -425 295 -421
rect 299 -425 303 -421
rect 328 -423 330 -421
rect 334 -423 336 -421
rect 51 -427 129 -425
rect 131 -427 135 -425
rect 256 -427 258 -425
rect 260 -427 309 -425
rect 315 -427 324 -425
rect 328 -427 340 -425
rect 354 -435 393 -124
rect 0 -448 393 -435
rect 0 -452 49 -448
rect 55 -452 102 -448
rect 0 -458 47 -452
rect 51 -458 53 -452
rect 57 -454 102 -452
rect 57 -458 68 -454
rect 72 -456 74 -454
rect 82 -456 94 -454
rect 100 -456 102 -454
rect 107 -454 180 -448
rect 197 -452 309 -448
rect 84 -458 92 -456
rect 0 -464 45 -458
rect 49 -462 55 -458
rect 59 -464 68 -458
rect 74 -460 80 -458
rect 0 -470 43 -464
rect 47 -470 57 -466
rect 61 -470 68 -464
rect 0 -472 41 -470
rect 45 -472 59 -470
rect 64 -472 68 -470
rect 72 -472 80 -460
rect 84 -468 90 -458
rect 96 -460 100 -458
rect 94 -466 102 -460
rect 96 -468 100 -466
rect 84 -470 92 -468
rect 84 -472 94 -470
rect 100 -472 102 -470
rect 107 -472 111 -454
rect 115 -456 117 -454
rect 123 -456 129 -454
rect 135 -456 141 -454
rect 123 -458 127 -456
rect 137 -458 141 -456
rect 145 -458 152 -454
rect 117 -460 125 -458
rect 129 -460 135 -458
rect 115 -468 125 -460
rect 139 -464 143 -458
rect 129 -466 143 -464
rect 148 -460 152 -458
rect 158 -458 164 -454
rect 168 -458 180 -454
rect 184 -454 309 -452
rect 184 -456 207 -454
rect 213 -456 221 -454
rect 225 -456 227 -454
rect 184 -458 205 -456
rect 215 -458 221 -456
rect 234 -458 236 -454
rect 240 -456 242 -454
rect 250 -456 258 -454
rect 268 -456 277 -454
rect 281 -456 283 -454
rect 291 -456 301 -454
rect 307 -456 309 -454
rect 313 -454 393 -448
rect 313 -456 324 -454
rect 330 -456 338 -454
rect 158 -460 162 -458
rect 148 -466 150 -460
rect 154 -466 156 -460
rect 160 -466 162 -460
rect 166 -466 180 -458
rect 195 -462 203 -458
rect 207 -460 213 -458
rect 131 -468 135 -466
rect 139 -468 145 -466
rect 115 -470 127 -468
rect 137 -470 145 -468
rect 115 -472 129 -470
rect 135 -472 145 -470
rect 152 -472 158 -466
rect 164 -472 180 -466
rect 184 -468 203 -462
rect 217 -464 221 -458
rect 227 -460 236 -458
rect 242 -460 248 -458
rect 207 -466 221 -464
rect 209 -468 213 -466
rect 217 -468 221 -466
rect 184 -470 205 -468
rect 215 -470 221 -468
rect 184 -472 207 -470
rect 213 -472 221 -470
rect 225 -472 236 -460
rect 240 -472 248 -460
rect 252 -460 256 -456
rect 260 -460 266 -458
rect 252 -462 262 -460
rect 252 -464 258 -462
rect 252 -470 256 -464
rect 262 -466 266 -464
rect 260 -468 266 -466
rect 270 -470 277 -456
rect 293 -458 299 -456
rect 313 -458 322 -456
rect 332 -458 338 -456
rect 352 -458 393 -454
rect 283 -460 289 -458
rect 252 -472 258 -470
rect 266 -472 268 -470
rect 272 -472 277 -470
rect 281 -472 289 -460
rect 293 -468 297 -458
rect 303 -460 307 -458
rect 301 -466 309 -460
rect 303 -468 307 -466
rect 313 -468 320 -458
rect 324 -460 330 -458
rect 334 -460 346 -458
rect 334 -462 344 -460
rect 350 -462 393 -458
rect 334 -464 342 -462
rect 348 -464 393 -462
rect 324 -466 340 -464
rect 346 -466 393 -464
rect 326 -468 330 -466
rect 334 -468 340 -466
rect 344 -468 393 -466
rect 293 -470 299 -468
rect 313 -470 322 -468
rect 332 -470 338 -468
rect 293 -472 301 -470
rect 307 -472 309 -470
rect 313 -472 324 -470
rect 330 -472 338 -470
rect 352 -472 393 -468
rect 0 -489 393 -472
rect 0 -513 84 -489
rect 102 -493 107 -489
rect 88 -499 107 -493
rect 102 -503 107 -499
rect 88 -509 107 -503
rect 102 -513 107 -509
rect 111 -493 117 -489
rect 121 -491 150 -489
rect 152 -491 176 -489
rect 188 -491 252 -489
rect 121 -493 148 -491
rect 111 -495 148 -493
rect 152 -495 172 -491
rect 191 -493 250 -491
rect 176 -495 186 -493
rect 193 -495 250 -493
rect 254 -495 393 -489
rect 111 -513 117 -495
rect 121 -497 131 -495
rect 139 -497 145 -495
rect 121 -499 129 -497
rect 141 -499 145 -497
rect 156 -499 170 -495
rect 176 -497 188 -495
rect 191 -497 201 -495
rect 207 -497 217 -495
rect 221 -497 223 -495
rect 229 -497 231 -495
rect 242 -497 248 -495
rect 121 -509 127 -499
rect 133 -501 137 -499
rect 131 -507 139 -501
rect 133 -509 137 -507
rect 143 -509 148 -499
rect 152 -507 170 -499
rect 174 -499 199 -497
rect 209 -499 217 -497
rect 244 -499 248 -497
rect 258 -499 260 -495
rect 264 -497 266 -495
rect 275 -497 287 -495
rect 293 -497 301 -495
rect 305 -497 307 -495
rect 277 -499 285 -497
rect 295 -499 301 -497
rect 313 -499 393 -495
rect 174 -501 197 -499
rect 201 -501 207 -499
rect 174 -505 182 -501
rect 176 -507 188 -505
rect 152 -509 172 -507
rect 176 -509 186 -507
rect 193 -509 197 -501
rect 211 -505 217 -499
rect 223 -501 229 -499
rect 234 -501 240 -499
rect 244 -501 250 -499
rect 201 -507 217 -505
rect 203 -509 207 -507
rect 211 -509 217 -507
rect 121 -511 129 -509
rect 141 -511 148 -509
rect 156 -511 172 -509
rect 193 -511 199 -509
rect 209 -511 217 -509
rect 121 -513 131 -511
rect 139 -513 150 -511
rect 156 -513 176 -511
rect 188 -513 201 -511
rect 207 -513 217 -511
rect 221 -503 229 -501
rect 238 -503 250 -501
rect 221 -505 231 -503
rect 242 -505 250 -503
rect 221 -507 238 -505
rect 221 -511 229 -507
rect 234 -509 240 -507
rect 244 -511 250 -505
rect 254 -509 260 -499
rect 266 -501 272 -499
rect 221 -513 231 -511
rect 242 -513 252 -511
rect 258 -513 260 -509
rect 264 -513 272 -501
rect 277 -509 283 -499
rect 287 -501 293 -499
rect 297 -505 301 -499
rect 307 -501 393 -499
rect 287 -507 301 -505
rect 289 -509 293 -507
rect 297 -509 301 -507
rect 277 -511 285 -509
rect 295 -511 301 -509
rect 277 -513 287 -511
rect 293 -513 301 -511
rect 305 -513 393 -501
rect 0 -544 393 -513
rect 0 -569 88 -544
rect 94 -548 104 -544
rect 92 -560 94 -552
rect 96 -554 102 -548
rect 111 -550 170 -544
rect 111 -552 119 -550
rect 129 -552 137 -550
rect 141 -552 143 -550
rect 150 -552 154 -550
rect 162 -552 170 -550
rect 174 -546 203 -544
rect 211 -546 242 -544
rect 250 -546 262 -544
rect 270 -546 281 -544
rect 289 -546 301 -544
rect 309 -546 393 -544
rect 174 -548 201 -546
rect 213 -548 240 -546
rect 252 -548 260 -546
rect 272 -548 279 -546
rect 291 -548 299 -546
rect 311 -548 393 -546
rect 174 -550 199 -548
rect 205 -550 211 -548
rect 174 -552 176 -550
rect 184 -552 199 -550
rect 203 -552 211 -550
rect 98 -560 100 -554
rect 104 -560 107 -552
rect 92 -566 96 -560
rect 102 -566 107 -560
rect 92 -569 98 -566
rect 100 -569 107 -566
rect 111 -556 117 -552
rect 121 -556 127 -554
rect 111 -558 123 -556
rect 111 -560 119 -558
rect 111 -566 117 -560
rect 123 -562 127 -560
rect 121 -564 127 -562
rect 131 -566 137 -552
rect 148 -554 152 -552
rect 143 -556 150 -554
rect 156 -556 160 -554
rect 164 -556 170 -552
rect 186 -554 211 -552
rect 215 -552 238 -548
rect 244 -550 250 -548
rect 242 -552 250 -550
rect 215 -554 250 -552
rect 254 -554 258 -548
rect 264 -550 268 -548
rect 176 -556 182 -554
rect 111 -569 119 -566
rect 127 -569 129 -566
rect 133 -569 137 -566
rect 141 -564 150 -556
rect 154 -562 170 -556
rect 156 -564 160 -562
rect 141 -566 152 -564
rect 164 -566 170 -562
rect 141 -569 154 -566
rect 162 -569 170 -566
rect 174 -569 182 -556
rect 186 -556 209 -554
rect 213 -556 248 -554
rect 186 -558 207 -556
rect 213 -558 246 -556
rect 252 -558 258 -554
rect 186 -560 205 -558
rect 211 -560 244 -558
rect 250 -560 258 -558
rect 186 -562 203 -560
rect 209 -562 242 -560
rect 248 -562 258 -560
rect 262 -562 270 -550
rect 186 -564 201 -562
rect 205 -564 240 -562
rect 244 -564 258 -562
rect 264 -564 268 -562
rect 275 -564 277 -548
rect 283 -550 287 -548
rect 281 -562 289 -550
rect 283 -564 287 -562
rect 293 -564 297 -548
rect 303 -550 307 -548
rect 301 -562 309 -550
rect 303 -564 307 -562
rect 313 -564 393 -548
rect 186 -569 199 -564
rect 215 -569 221 -564
rect 225 -569 238 -564
rect 254 -566 260 -564
rect 272 -566 279 -564
rect 291 -566 299 -564
rect 311 -566 393 -564
rect 254 -569 262 -566
rect 270 -569 281 -566
rect 289 -569 301 -566
rect 309 -569 393 -566
rect 0 -571 223 -569
rect 0 -575 221 -571
rect 225 -573 393 -569
rect 223 -575 393 -573
rect 0 -587 393 -575
<< end >>
