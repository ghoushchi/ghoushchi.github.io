magic
tech scmos
timestamp 951985653
<< metal1 >>
rect 1732 2927 1755 2933
rect 1732 2925 1758 2927
rect 361 2909 365 2915
rect 802 2912 805 2915
rect 995 2912 998 2915
rect 1372 2912 1375 2915
rect 347 2905 365 2909
rect 1749 2909 1758 2925
rect 1942 2912 1945 2915
rect 2135 2912 2138 2915
rect 2512 2912 2515 2915
rect 2705 2912 2708 2915
rect 1618 2791 1666 2900
rect 320 2645 335 2649
rect 835 2639 839 2652
rect 875 2632 879 2644
rect 963 2639 967 2676
rect 987 2639 991 2668
rect 1051 2636 1055 2660
rect 1075 2639 1079 2684
rect 1139 2638 1143 2692
rect 1163 2638 1167 2700
rect 1251 2639 1255 2708
rect 1259 2637 1263 2716
rect 1267 2638 1271 2724
rect 1275 2639 1279 2732
rect 1283 2636 1287 2740
rect 1299 2636 1303 2748
rect 1307 2639 1311 2756
rect 1315 2636 1319 2764
rect 571 2601 759 2606
rect 773 2601 775 2606
rect 571 2596 775 2601
rect 779 2597 805 2606
rect 779 2596 801 2597
rect 1618 2593 1666 2772
rect 1725 2815 1745 2900
rect 1745 2795 1930 2815
rect 1937 2795 2051 2815
rect 2057 2795 2171 2815
rect 2177 2795 2291 2815
rect 2297 2795 2411 2815
rect 2417 2795 2561 2815
rect 2567 2795 2603 2815
rect 1725 2606 1745 2795
rect 1779 2772 1992 2791
rect 1997 2772 2111 2791
rect 2117 2772 2231 2791
rect 2237 2772 2351 2791
rect 2357 2772 2470 2791
rect 2476 2772 2582 2791
rect 1914 2764 2449 2768
rect 1914 2756 2377 2760
rect 1914 2748 2329 2752
rect 1914 2740 2257 2744
rect 1914 2732 2209 2736
rect 1914 2724 2137 2728
rect 1913 2716 2089 2720
rect 1913 2708 2017 2712
rect 1913 2700 2545 2704
rect 1913 2692 2537 2696
rect 1913 2684 2529 2688
rect 1912 2676 2521 2680
rect 1913 2668 2513 2672
rect 1912 2660 2505 2664
rect 1913 2652 2497 2656
rect 1912 2644 2489 2648
rect 1912 2636 2481 2640
rect 1745 2597 1810 2606
rect 320 2581 327 2585
rect 595 2582 693 2592
rect 347 2574 578 2578
rect 1666 2575 1752 2593
rect 1758 2575 1872 2593
rect 1549 2566 1915 2570
rect 339 2542 578 2546
rect 331 2510 573 2514
rect 1549 2510 1907 2514
rect 331 2478 576 2482
rect 339 2446 657 2450
rect 1549 2446 1840 2450
rect 1637 2423 1725 2443
rect 347 2414 574 2418
rect 355 2382 573 2386
rect 363 2350 574 2354
rect 320 2076 327 2080
rect 320 2010 335 2014
rect 1530 1803 1617 1809
rect 1530 1792 1592 1799
rect 1529 1692 1592 1698
rect 1228 1630 1236 1634
rect 1240 1630 1362 1634
rect 1366 1630 1504 1634
rect 1228 1622 1274 1626
rect 1278 1622 1370 1626
rect 1374 1622 1504 1626
rect 1655 1620 1663 1624
rect 1228 1614 1312 1618
rect 1316 1614 1378 1618
rect 1382 1614 1504 1618
rect 1228 1606 1350 1610
rect 1354 1606 1504 1610
rect 1228 1598 1388 1602
rect 1392 1598 1503 1602
rect 1539 1599 1592 1618
rect 1228 1590 1427 1594
rect 1431 1590 1504 1594
rect 1647 1588 1663 1592
rect 1228 1582 1467 1586
rect 1471 1582 1504 1586
rect 1228 1574 1499 1578
rect 1503 1574 1504 1578
rect 607 1567 675 1571
rect 991 1566 1066 1570
rect 1095 1566 1185 1570
rect 1197 1566 1306 1570
rect 1414 1566 1467 1570
rect 1565 1566 1617 1587
rect 623 1557 705 1561
rect 727 1557 762 1561
rect 911 1558 936 1562
rect 951 1558 994 1562
rect 1055 1558 1114 1562
rect 1159 1558 1234 1562
rect 1351 1560 1386 1564
rect 1422 1559 1499 1563
rect 733 1549 739 1553
rect 754 1548 849 1553
rect 855 1548 969 1553
rect 975 1548 1089 1553
rect 1095 1548 1209 1553
rect 1215 1548 1329 1553
rect 1334 1548 1519 1553
rect 742 1539 749 1544
rect 795 1541 800 1545
rect 810 1541 909 1545
rect 795 1540 909 1541
rect 915 1540 1029 1545
rect 1035 1540 1149 1545
rect 1155 1541 1201 1545
rect 1205 1541 1269 1545
rect 1155 1540 1269 1541
rect 1275 1540 1545 1545
rect 671 1533 713 1537
rect 1435 1530 1659 1534
rect 1443 1522 1651 1526
rect 1451 1514 1643 1518
rect 320 1505 343 1509
rect 320 1440 351 1444
rect 695 1303 724 1307
rect 687 1207 724 1211
rect 1362 1087 1418 1091
rect 1363 1079 1410 1083
rect 1364 1071 1402 1075
rect 2888 1073 2905 1076
rect 1363 1063 1394 1067
rect 1581 1060 1660 1064
rect 1799 1060 1907 1064
rect 1362 1055 1386 1059
rect 1589 1052 1659 1056
rect 1363 1047 1378 1051
rect 1597 1044 1659 1048
rect 1362 1039 1370 1043
rect 1605 1036 1659 1040
rect 709 1023 724 1027
rect 1358 1023 1431 1027
rect 717 1015 724 1019
rect 1350 1015 1439 1019
rect 1342 1008 1447 1012
rect 1399 1000 1674 1004
rect 1407 992 1682 996
rect 1573 984 1666 988
rect 320 935 359 939
rect 1613 916 1659 920
rect 1621 900 1659 904
rect 320 870 327 874
rect 575 863 595 891
rect 1629 884 1659 888
rect 1637 868 1660 872
rect 568 851 595 863
rect 1645 852 1659 856
rect 568 843 724 851
rect 1364 843 1519 848
rect 592 839 724 840
rect 592 831 732 839
rect 1376 836 1742 840
rect 766 828 1372 832
rect 1384 828 1734 832
rect 1904 825 1916 828
rect 331 821 729 825
rect 733 821 1130 825
rect 1134 821 1380 825
rect 1904 824 1907 825
rect 1911 824 1914 825
rect 537 813 1066 817
rect 703 805 770 809
rect 926 805 1020 809
rect 1350 808 1519 817
rect 1539 808 1899 817
rect 647 794 675 798
rect 1364 795 1545 804
rect 1565 795 1883 804
rect 331 786 755 790
rect 759 786 762 790
rect 733 772 763 776
rect 1047 773 1170 777
rect 1104 763 1114 767
rect 529 755 644 759
rect 1503 739 1601 743
rect 1503 731 1577 735
rect 2896 734 2905 737
rect 592 717 601 721
rect 1504 717 1545 721
rect 1659 700 1703 709
rect 1817 700 1818 709
rect 2566 700 2603 709
rect 568 665 597 669
rect 1504 665 1519 669
rect 1660 667 1757 676
rect 2476 667 2582 676
rect 1503 651 1569 655
rect 2456 649 2884 653
rect 1503 643 1585 647
rect 2376 640 2892 644
rect 1503 635 1593 639
rect 2336 631 2892 635
rect 1503 627 1617 631
rect 1503 619 1609 623
rect 1503 611 1633 615
rect 592 597 596 601
rect 1504 597 1545 601
rect 568 545 596 549
rect 1504 545 1519 549
rect 1503 531 1641 535
rect 1503 523 1734 526
rect 1502 515 1625 519
rect 2896 503 2905 506
rect 2896 502 2899 503
rect 537 498 699 502
rect 529 491 1068 495
rect 1400 493 1863 496
rect 1392 486 1855 489
rect 592 465 1545 483
rect 1565 465 1580 483
rect 1628 465 1805 483
rect 1827 465 2603 483
rect 568 442 1473 460
rect 1485 442 1519 460
rect 1539 442 1777 460
rect 1800 442 2581 460
rect 320 365 327 369
rect 1299 340 2009 345
rect 361 329 699 333
rect 361 320 364 329
rect 729 319 732 328
rect 1068 319 1071 325
rect 1299 319 1302 340
rect 2253 338 2782 342
rect 1473 250 1485 327
rect 1869 328 2089 333
rect 2133 330 2211 334
rect 2221 330 2442 334
rect 1869 319 1872 328
rect 2208 320 2211 330
rect 2439 315 2442 330
rect 2778 319 2782 338
<< metal2 >>
rect 446 3134 500 3187
rect 1580 3134 1634 3187
rect 424 2981 428 2985
rect 801 2912 805 2915
rect 994 2912 998 2915
rect 1371 2912 1375 2915
rect 1618 2909 1666 2915
rect 1941 2912 1945 2915
rect 49 2744 103 2797
rect 250 2709 254 2713
rect 250 2517 254 2521
rect 327 2514 331 2581
rect 335 2546 339 2645
rect 343 2578 347 2905
rect 1745 2900 1749 2909
rect 2134 2912 2138 2915
rect 2511 2912 2515 2915
rect 2704 2912 2708 2915
rect 1666 2772 1770 2791
rect 1319 2764 1910 2768
rect 1311 2756 1910 2760
rect 1303 2748 1910 2752
rect 1287 2740 1910 2744
rect 1279 2732 1910 2736
rect 1271 2724 1910 2728
rect 1263 2716 1909 2720
rect 1255 2708 1909 2712
rect 1167 2700 1909 2704
rect 1143 2692 1909 2696
rect 1079 2684 1909 2688
rect 967 2676 1908 2680
rect 991 2668 1909 2672
rect 1055 2660 1908 2664
rect 839 2652 1909 2656
rect 879 2644 1908 2648
rect 903 2636 1908 2640
rect 773 2601 786 2606
rect 817 2597 1725 2606
rect 54 2453 108 2506
rect 54 2166 108 2219
rect 250 2139 254 2143
rect 327 2080 331 2478
rect 335 2014 339 2446
rect 250 1947 254 1951
rect 63 1875 117 1928
rect 51 1597 105 1650
rect 250 1569 254 1573
rect 343 1509 347 2414
rect 351 1444 355 2382
rect 250 1377 254 1381
rect 57 1307 111 1360
rect 48 1020 102 1073
rect 250 999 254 1003
rect 359 939 363 2350
rect 551 1809 571 2596
rect 703 2582 706 2592
rect 1245 2582 1618 2593
rect 551 1803 560 1809
rect 575 1800 595 2582
rect 1245 2581 1436 2582
rect 1592 2575 1618 2582
rect 586 1794 595 1800
rect 1592 1799 1613 2575
rect 1725 2443 1745 2597
rect 1592 1698 1613 1792
rect 551 1628 569 1631
rect 551 887 571 1628
rect 575 911 595 1580
rect 619 1561 623 1568
rect 667 1537 671 1568
rect 327 825 331 870
rect 551 867 592 887
rect 250 807 254 811
rect 45 735 99 788
rect 50 452 104 505
rect 250 429 254 433
rect 327 369 331 786
rect 525 495 529 755
rect 533 502 537 813
rect 548 669 568 843
rect 548 549 568 665
rect 548 460 568 545
rect 572 840 592 867
rect 572 721 592 831
rect 675 798 679 1567
rect 643 766 647 794
rect 683 790 687 1207
rect 676 786 687 790
rect 676 766 680 786
rect 691 782 695 1303
rect 705 1027 709 1557
rect 715 1545 719 1568
rect 723 1561 727 1568
rect 739 1553 743 1568
rect 749 1553 754 1580
rect 715 1541 725 1545
rect 713 1019 717 1533
rect 721 1011 725 1541
rect 729 825 733 1549
rect 749 1544 754 1548
rect 737 1414 742 1539
rect 762 1421 766 1557
rect 800 1545 810 1693
rect 827 1545 831 1568
rect 849 1540 855 1548
rect 859 1549 863 1568
rect 907 1562 911 1568
rect 947 1562 951 1568
rect 1051 1562 1055 1569
rect 859 1545 878 1549
rect 936 1545 940 1558
rect 872 1544 876 1545
rect 936 1541 947 1545
rect 969 1540 975 1548
rect 994 1545 998 1558
rect 1066 1545 1070 1566
rect 1155 1562 1159 1568
rect 1089 1540 1095 1548
rect 1114 1545 1118 1558
rect 1185 1545 1189 1566
rect 1201 1545 1205 1693
rect 1209 1540 1215 1548
rect 1234 1545 1238 1558
rect 1306 1545 1310 1566
rect 1329 1553 1334 1692
rect 1347 1564 1351 1569
rect 1329 1540 1334 1548
rect 1362 1035 1366 1630
rect 1362 1026 1366 1031
rect 1370 1043 1374 1622
rect 1592 1618 1613 1692
rect 1370 1026 1374 1039
rect 1378 1051 1382 1614
rect 1617 1809 1637 2423
rect 1402 1574 1431 1578
rect 1387 1568 1398 1572
rect 1378 1026 1382 1047
rect 1386 1059 1390 1560
rect 1386 1026 1390 1055
rect 1394 1067 1398 1568
rect 1394 1026 1398 1063
rect 1402 1075 1406 1574
rect 1402 1026 1406 1071
rect 1410 1083 1414 1566
rect 1499 1563 1503 1568
rect 1410 1026 1414 1079
rect 1418 1091 1422 1559
rect 1519 1553 1539 1598
rect 1617 1587 1637 1803
rect 1418 1026 1422 1087
rect 1431 1027 1435 1530
rect 1439 1019 1443 1522
rect 1447 1012 1451 1514
rect 1130 927 1134 994
rect 1114 923 1134 927
rect 684 778 695 782
rect 684 766 688 778
rect 699 766 703 805
rect 729 776 733 821
rect 762 790 766 828
rect 770 809 774 825
rect 802 809 806 825
rect 796 805 806 809
rect 759 786 762 790
rect 755 765 759 786
rect 763 766 767 772
rect 796 766 800 805
rect 810 801 814 825
rect 922 809 926 825
rect 1066 817 1070 825
rect 804 797 814 801
rect 804 766 808 797
rect 1020 770 1024 805
rect 1020 763 1023 770
rect 1043 766 1047 773
rect 1114 767 1118 923
rect 1130 825 1134 887
rect 1170 777 1174 825
rect 1341 817 1350 843
rect 1355 804 1364 835
rect 1372 832 1376 836
rect 1380 825 1384 828
rect 1395 766 1399 1000
rect 1403 766 1407 992
rect 1519 848 1539 1548
rect 1519 817 1539 843
rect 572 601 592 717
rect 572 483 592 597
rect 1519 669 1539 808
rect 1519 549 1539 665
rect 699 333 703 498
rect 795 332 799 499
rect 733 328 799 332
rect 1068 329 1072 491
rect 1388 490 1391 499
rect 1396 497 1399 499
rect 1519 460 1539 545
rect 1545 1545 1565 1566
rect 1545 804 1565 1540
rect 1643 1518 1647 1588
rect 1651 1526 1655 1620
rect 1659 1534 1663 1668
rect 1752 1429 1758 2575
rect 1810 1428 1818 2597
rect 1840 1706 1844 2446
rect 1872 1879 1878 2575
rect 1907 2156 1911 2510
rect 1915 2336 1919 2566
rect 1930 2454 1937 2795
rect 1992 2630 1997 2772
rect 2017 2636 2021 2708
rect 2051 2630 2057 2795
rect 2089 2636 2093 2716
rect 2111 2630 2117 2772
rect 2137 2636 2141 2724
rect 2171 2630 2177 2795
rect 2209 2636 2213 2732
rect 2231 2630 2237 2772
rect 2257 2636 2261 2740
rect 2291 2630 2297 2795
rect 2329 2636 2333 2748
rect 2351 2630 2357 2772
rect 2377 2636 2381 2756
rect 2411 2630 2417 2795
rect 2449 2636 2453 2764
rect 2470 2629 2476 2772
rect 2481 2632 2485 2636
rect 2489 2631 2493 2644
rect 2497 2633 2501 2652
rect 2505 2633 2509 2660
rect 2513 2634 2517 2668
rect 2521 2635 2525 2676
rect 2529 2636 2533 2684
rect 2537 2636 2541 2692
rect 2545 2636 2549 2700
rect 2561 2600 2566 2795
rect 1545 721 1565 795
rect 1545 601 1565 717
rect 1569 655 1573 984
rect 1577 735 1581 1060
rect 1585 647 1589 1052
rect 1593 639 1597 1044
rect 1601 743 1605 1036
rect 1666 988 1670 1016
rect 1609 623 1613 916
rect 1617 631 1621 900
rect 1545 483 1565 597
rect 1625 519 1629 884
rect 1633 615 1637 868
rect 1641 535 1645 852
rect 1734 697 1738 828
rect 1742 690 1746 836
rect 1907 825 1911 1060
rect 1810 700 1818 709
rect 1734 527 1738 679
rect 1805 671 1811 700
rect 1473 336 1485 442
rect 1580 320 1628 465
rect 1777 460 1800 667
rect 1817 662 1827 700
rect 1805 483 1827 662
rect 1855 490 1859 788
rect 1863 497 1867 748
rect 1883 709 1892 795
rect 1899 676 1908 808
rect 2582 676 2599 2772
rect 2009 345 2013 666
rect 2089 333 2093 666
rect 2129 334 2133 666
rect 2209 334 2213 665
rect 2249 342 2253 664
rect 2332 635 2336 662
rect 2372 644 2376 662
rect 2452 653 2456 662
rect 2582 460 2599 667
rect 2603 709 2621 2795
rect 2971 2709 2975 2713
rect 2971 2517 2975 2521
rect 2971 2139 2975 2143
rect 2971 1947 2975 1951
rect 2971 1569 2975 1573
rect 2971 1377 2975 1381
rect 2603 483 2621 700
rect 2884 653 2888 1072
rect 3124 1028 3178 1081
rect 2963 999 2967 1003
rect 2963 807 2967 811
rect 3125 741 3179 794
rect 2892 644 2896 733
rect 2892 506 2896 631
rect 3125 460 3179 513
rect 2963 429 2967 433
rect 2209 330 2217 334
rect 424 314 429 320
rect 802 258 807 262
rect 994 258 998 262
rect 1372 258 1376 262
rect 1942 258 1946 262
rect 2134 258 2138 262
rect 2512 258 2516 262
rect 2704 258 2708 262
rect 424 250 428 254
rect 450 44 504 97
rect 732 48 786 101
rect 1022 46 1076 99
rect 1306 51 1360 104
rect 1589 48 1643 101
rect 1869 53 1923 106
rect 2149 58 2203 111
rect 2448 54 2502 107
rect 2732 52 2786 105
<< m2contact >>
rect 343 2905 347 2909
rect 801 2908 805 2912
rect 994 2908 998 2912
rect 1371 2908 1375 2912
rect 1618 2900 1666 2909
rect 1618 2772 1666 2791
rect 1315 2764 1319 2768
rect 1307 2756 1311 2760
rect 1299 2748 1303 2752
rect 1283 2740 1287 2744
rect 1275 2732 1279 2736
rect 1267 2724 1271 2728
rect 1259 2716 1263 2720
rect 1251 2708 1255 2712
rect 1163 2700 1167 2704
rect 1139 2692 1143 2696
rect 1075 2684 1079 2688
rect 963 2676 967 2680
rect 835 2652 839 2656
rect 335 2645 339 2649
rect 875 2644 879 2648
rect 899 2636 903 2640
rect 987 2668 991 2672
rect 1051 2660 1055 2664
rect 551 2596 571 2606
rect 759 2601 773 2606
rect 805 2597 817 2606
rect 1725 2900 1745 2909
rect 1749 2900 1758 2909
rect 1941 2908 1945 2912
rect 2134 2908 2138 2912
rect 2511 2908 2515 2912
rect 2704 2908 2708 2912
rect 1725 2795 1745 2815
rect 1930 2795 1937 2815
rect 2051 2795 2057 2815
rect 2171 2795 2177 2815
rect 2291 2795 2297 2815
rect 2411 2795 2417 2815
rect 2561 2795 2567 2815
rect 2603 2795 2621 2815
rect 1770 2772 1779 2791
rect 1992 2772 1997 2791
rect 2111 2772 2117 2791
rect 2231 2772 2237 2791
rect 2351 2772 2357 2791
rect 2470 2772 2476 2791
rect 2582 2772 2599 2791
rect 1910 2764 1914 2768
rect 2449 2764 2453 2768
rect 1910 2756 1914 2760
rect 2377 2756 2381 2760
rect 1910 2748 1914 2752
rect 2329 2748 2333 2752
rect 1910 2740 1914 2744
rect 2257 2740 2261 2744
rect 1910 2732 1914 2736
rect 2209 2732 2213 2736
rect 1910 2724 1914 2728
rect 2137 2724 2141 2728
rect 1909 2716 1913 2720
rect 2089 2716 2093 2720
rect 1909 2708 1913 2712
rect 2017 2708 2021 2712
rect 1909 2700 1913 2704
rect 2545 2700 2549 2704
rect 1909 2692 1913 2696
rect 2537 2692 2541 2696
rect 1909 2684 1913 2688
rect 2529 2684 2533 2688
rect 1908 2676 1912 2680
rect 2521 2676 2525 2680
rect 1909 2668 1913 2672
rect 2513 2668 2517 2672
rect 1908 2660 1912 2664
rect 2505 2660 2509 2664
rect 1909 2652 1913 2656
rect 2497 2652 2501 2656
rect 1908 2644 1912 2648
rect 2489 2644 2493 2648
rect 1908 2636 1912 2640
rect 2481 2636 2485 2640
rect 1725 2597 1745 2606
rect 1810 2597 1818 2606
rect 327 2581 331 2585
rect 575 2582 595 2592
rect 693 2582 703 2592
rect 343 2574 347 2578
rect 1618 2575 1666 2593
rect 1752 2575 1758 2593
rect 1872 2575 1878 2593
rect 1545 2566 1549 2570
rect 1915 2566 1919 2570
rect 335 2542 339 2546
rect 327 2510 331 2514
rect 1545 2510 1549 2514
rect 1907 2510 1911 2514
rect 327 2478 331 2482
rect 335 2446 339 2450
rect 1545 2446 1549 2450
rect 1840 2446 1844 2450
rect 1617 2423 1637 2443
rect 1725 2423 1745 2443
rect 343 2414 347 2418
rect 351 2382 355 2386
rect 359 2350 363 2354
rect 1915 2332 1919 2336
rect 1907 2152 1911 2156
rect 327 2076 331 2080
rect 335 2010 339 2014
rect 1524 1803 1530 1809
rect 1617 1803 1637 1809
rect 1524 1792 1530 1799
rect 1592 1792 1613 1799
rect 1840 1702 1844 1706
rect 1329 1692 1334 1696
rect 1592 1692 1613 1698
rect 1659 1668 1663 1672
rect 1236 1630 1240 1634
rect 1362 1630 1366 1634
rect 1274 1622 1278 1626
rect 1370 1622 1374 1626
rect 1651 1620 1655 1624
rect 1312 1614 1316 1618
rect 1378 1614 1382 1618
rect 1350 1606 1354 1610
rect 1388 1598 1392 1602
rect 1519 1598 1539 1618
rect 1592 1599 1613 1618
rect 1427 1590 1431 1594
rect 1643 1588 1647 1592
rect 749 1580 754 1585
rect 1467 1582 1471 1586
rect 1499 1574 1503 1578
rect 603 1567 607 1571
rect 675 1567 679 1571
rect 987 1566 991 1570
rect 1066 1566 1070 1570
rect 1091 1566 1095 1570
rect 1185 1566 1189 1570
rect 1193 1566 1197 1570
rect 1306 1566 1310 1570
rect 1410 1566 1414 1570
rect 1467 1566 1471 1570
rect 1545 1566 1565 1587
rect 1617 1566 1637 1587
rect 619 1557 623 1561
rect 705 1557 709 1561
rect 723 1557 727 1561
rect 762 1557 766 1561
rect 907 1558 911 1562
rect 936 1558 940 1562
rect 947 1558 951 1562
rect 994 1558 998 1562
rect 1051 1558 1055 1562
rect 1114 1558 1118 1562
rect 1155 1558 1159 1562
rect 1234 1558 1238 1562
rect 1347 1560 1351 1564
rect 1386 1560 1390 1564
rect 1418 1559 1422 1563
rect 1499 1559 1503 1563
rect 729 1549 733 1553
rect 739 1549 743 1553
rect 749 1548 754 1553
rect 849 1548 855 1553
rect 969 1548 975 1553
rect 1089 1548 1095 1553
rect 1209 1548 1215 1553
rect 1329 1548 1334 1553
rect 1519 1548 1539 1553
rect 737 1539 742 1544
rect 749 1539 754 1544
rect 790 1540 795 1545
rect 800 1541 810 1545
rect 909 1540 915 1545
rect 1029 1540 1035 1545
rect 1149 1540 1155 1545
rect 1201 1541 1205 1545
rect 1269 1540 1275 1545
rect 1545 1540 1565 1545
rect 667 1533 671 1537
rect 713 1533 717 1537
rect 1431 1530 1435 1534
rect 1659 1530 1663 1534
rect 1439 1522 1443 1526
rect 1651 1522 1655 1526
rect 1447 1514 1451 1518
rect 1643 1514 1647 1518
rect 343 1505 347 1509
rect 351 1440 355 1444
rect 691 1303 695 1307
rect 683 1207 687 1211
rect 1418 1087 1422 1091
rect 1410 1079 1414 1083
rect 1402 1071 1406 1075
rect 2884 1072 2888 1076
rect 1394 1063 1398 1067
rect 1577 1060 1581 1064
rect 1907 1060 1911 1064
rect 1386 1055 1390 1059
rect 1585 1052 1589 1056
rect 1378 1047 1382 1051
rect 1593 1044 1597 1048
rect 1370 1039 1374 1043
rect 1601 1036 1605 1040
rect 1362 1031 1366 1035
rect 705 1023 709 1027
rect 1431 1023 1435 1027
rect 713 1015 717 1019
rect 1439 1015 1443 1019
rect 721 1007 725 1011
rect 1447 1008 1451 1012
rect 1395 1000 1399 1004
rect 1674 1000 1678 1004
rect 1403 992 1407 996
rect 1682 992 1686 996
rect 1569 984 1573 988
rect 1666 984 1670 988
rect 359 935 363 939
rect 1609 916 1613 920
rect 575 891 595 911
rect 1617 900 1621 904
rect 327 870 331 874
rect 1625 884 1629 888
rect 1633 868 1637 872
rect 548 843 568 863
rect 1641 852 1645 856
rect 1341 843 1350 848
rect 1519 843 1539 848
rect 572 831 592 840
rect 1355 835 1364 840
rect 1372 836 1376 840
rect 1742 836 1746 840
rect 762 828 766 832
rect 1372 828 1376 832
rect 1380 828 1384 832
rect 1734 828 1738 832
rect 327 821 331 825
rect 729 821 733 825
rect 1130 821 1134 825
rect 1380 821 1384 825
rect 1907 821 1911 825
rect 533 813 537 817
rect 1066 813 1070 817
rect 699 805 703 809
rect 770 805 774 809
rect 922 805 926 809
rect 1020 805 1024 809
rect 1341 808 1350 817
rect 1519 808 1539 817
rect 1899 808 1908 817
rect 643 794 647 798
rect 675 794 679 798
rect 1355 795 1364 804
rect 1545 795 1565 804
rect 1883 795 1892 804
rect 327 786 331 790
rect 755 786 759 790
rect 762 786 766 790
rect 1855 788 1859 792
rect 729 772 733 776
rect 763 772 767 776
rect 1043 773 1047 777
rect 1170 773 1174 777
rect 1114 763 1118 767
rect 525 755 529 759
rect 1863 748 1867 752
rect 1601 739 1605 743
rect 1577 731 1581 735
rect 2892 733 2896 737
rect 572 717 592 721
rect 1545 717 1565 721
rect 1805 700 1810 709
rect 1818 700 1827 709
rect 1883 700 1892 709
rect 2603 700 2621 709
rect 1734 693 1738 697
rect 1742 686 1746 690
rect 1734 679 1738 683
rect 548 665 568 669
rect 1519 665 1539 669
rect 1777 667 1800 676
rect 1899 667 1908 676
rect 2582 667 2599 676
rect 1569 651 1573 655
rect 2452 649 2456 653
rect 2884 649 2888 653
rect 1585 643 1589 647
rect 2372 640 2376 644
rect 2892 640 2896 644
rect 1593 635 1597 639
rect 2332 631 2336 635
rect 2892 631 2896 635
rect 1617 627 1621 631
rect 1609 619 1613 623
rect 1633 611 1637 615
rect 572 597 592 601
rect 1545 597 1565 601
rect 548 545 568 549
rect 1519 545 1539 549
rect 1641 531 1645 535
rect 1734 523 1738 527
rect 1625 515 1629 519
rect 2892 502 2896 506
rect 533 498 537 502
rect 699 498 703 502
rect 525 491 529 495
rect 1068 491 1072 495
rect 1396 493 1400 497
rect 1863 493 1867 497
rect 1388 486 1392 490
rect 1855 486 1859 490
rect 572 465 592 483
rect 1545 465 1565 483
rect 1580 465 1628 483
rect 1805 465 1827 483
rect 2603 465 2621 483
rect 548 442 568 460
rect 1473 442 1485 460
rect 1519 442 1539 460
rect 1777 442 1800 460
rect 2581 442 2599 460
rect 327 365 331 369
rect 2009 340 2014 345
rect 699 329 703 333
rect 729 328 733 332
rect 1068 325 1072 329
rect 2249 338 2253 342
rect 1473 327 1485 336
rect 2089 328 2093 333
rect 2128 330 2133 334
rect 2217 330 2221 334
rect 1473 244 1485 250
use tl 2_0
timestamp 950486748
transform 1 0 0 0 1 2900
box 0 0 330 335
use io 3_0
timestamp 950486748
transform 1 0 330 0 1 2915
box 0 0 285 320
use io 3_1
timestamp 950486748
transform -1 0 900 0 1 2915
box 0 0 285 320
use io 3_2
timestamp 950486748
transform 1 0 900 0 1 2915
box 0 0 285 320
use io 3_3
timestamp 950486748
transform -1 0 1470 0 1 2915
box 0 0 285 320
use gnd 4_0
timestamp 950486748
transform 1 0 1470 0 1 2915
box 0 0 285 320
use io 3_4
timestamp 950486748
transform -1 0 2040 0 1 2915
box 0 0 285 320
use io 3_5
timestamp 950486748
transform 1 0 2040 0 1 2915
box 0 0 285 320
use io 3_6
timestamp 950486748
transform -1 0 2610 0 1 2915
box 0 0 285 320
use io 3_7
timestamp 950486748
transform 1 0 2610 0 1 2915
box 0 0 285 320
use tr 5_0
timestamp 950486748
transform 1 0 2895 0 1 2900
box 0 0 330 335
use io 3_8
timestamp 950486748
transform 0 -1 320 1 0 2615
box 0 0 285 320
use io 3_9
timestamp 950486748
transform 0 -1 320 -1 0 2615
box 0 0 285 320
use io 3_10
timestamp 950486748
transform 0 -1 320 1 0 2045
box 0 0 285 320
use io 3_11
timestamp 950486748
transform 0 -1 320 -1 0 2045
box 0 0 285 320
use io 3_12
timestamp 950486748
transform 0 -1 320 1 0 1475
box 0 0 285 320
use art art_0
timestamp 951963504
transform 1 0 1443 0 1 2408
box 0 -587 393 2
use supremeMEM supremeMEM_0
timestamp 951985653
transform 1 0 573 0 1 1568
box -22 0 976 1072
use io 3_13
timestamp 950486748
transform 0 -1 320 -1 0 1475
box 0 0 285 320
use io 3_14
timestamp 950486748
transform 0 -1 320 1 0 905
box 0 0 285 320
use io 3_15
timestamp 950486748
transform 0 -1 320 -1 0 905
box 0 0 285 320
use counters counters_0
timestamp 951985653
transform 1 0 724 0 1 825
box 0 0 640 720
use io 3_16
timestamp 950486748
transform 0 -1 320 1 0 335
box 0 0 285 320
use controller controller_0
timestamp 951733675
transform 1 0 598 0 1 501
box -4 -2 906 266
use supremeDP supremeDP_0
timestamp 951985653
transform 0 -1 2571 -1 0 2638
box 0 0 1976 912
use io 3_17
timestamp 950486748
transform 0 1 2905 1 0 2615
box 0 0 285 320
use io 3_18
timestamp 950486748
transform 0 1 2905 -1 0 2615
box 0 0 285 320
use io 3_19
timestamp 950486748
transform 0 1 2905 1 0 2045
box 0 0 285 320
use io 3_20
timestamp 950486748
transform 0 1 2905 -1 0 2045
box 0 0 285 320
use io 3_21
timestamp 950486748
transform 0 1 2905 1 0 1475
box 0 0 285 320
use io 3_22
timestamp 950486748
transform 0 1 2905 -1 0 1475
box 0 0 285 320
use io 3_23
timestamp 950486748
transform 0 1 2905 1 0 905
box 0 0 285 320
use io 3_24
timestamp 950486748
transform 0 1 2905 -1 0 905
box 0 0 285 320
use io 3_25
timestamp 950486748
transform 0 1 2905 1 0 335
box 0 0 285 320
use bl 6_0
timestamp 950486748
transform 1 0 0 0 1 0
box 0 0 330 335
use io 3_26
timestamp 950486748
transform 1 0 330 0 -1 320
box 0 0 285 320
use io 3_27
timestamp 950486748
transform -1 0 900 0 -1 320
box 0 0 285 320
use io 3_28
timestamp 950486748
transform 1 0 900 0 -1 320
box 0 0 285 320
use io 3_29
timestamp 950486748
transform -1 0 1470 0 -1 320
box 0 0 285 320
use vdd 7_0
timestamp 950486748
transform 1 0 1470 0 -1 320
box 0 0 285 320
use io 3_30
timestamp 950486748
transform -1 0 2040 0 -1 320
box 0 0 285 320
use io 3_31
timestamp 950486748
transform 1 0 2040 0 -1 320
box 0 0 285 320
use io 3_32
timestamp 950486748
transform -1 0 2610 0 -1 320
box 0 0 285 320
use io 3_33
timestamp 950486748
transform 1 0 2610 0 -1 320
box 0 0 285 320
use br 8_0
timestamp 950486748
transform 1 0 2895 0 1 0
box 0 0 330 335
<< labels >>
rlabel metal2 1580 3134 1634 3187 0 Gnd
rlabel metal2 45 735 99 788 0 Phi1
rlabel metal2 50 452 104 505 0 Phi2
rlabel metal2 450 44 504 97 0 Reset_s1
rlabel metal2 732 48 786 101 0 Input_Ready_s1
rlabel metal2 1022 46 1076 99 0 Output_Ready_q1
rlabel metal2 1589 48 1643 101 0 Vdd
rlabel metal2 1306 51 1360 104 0 Final_Output_s1[7]
rlabel metal2 1869 53 1923 106 0 Final_Output_s1[6]
rlabel metal2 2149 58 2203 111 0 Final_Output_s1[5]
rlabel metal2 2448 54 2502 107 0 Final_Output_s1[4]
rlabel metal2 2732 52 2786 105 0 Final_Output_s1[3]
rlabel metal2 3125 460 3179 513 0 Final_Output_s1[2]
rlabel metal2 3125 741 3179 794 0 Final_Output_s1[1]
rlabel metal2 3124 1028 3178 1081 0 Final_Output_s1[0]
rlabel metal2 446 3134 500 3187 0 Pixel_s1[7]
rlabel metal2 49 2744 103 2797 0 Pixel_s1[6]
rlabel metal2 54 2453 108 2506 0 Pixel_s1[5]
rlabel metal2 54 2166 108 2219 0 Pixel_s1[4]
rlabel metal2 63 1875 117 1928 0 Pixel_s1[3]
rlabel metal2 51 1597 105 1650 0 Pixel_s1[2]
rlabel metal2 57 1307 111 1360 0 Pixel_s1[1]
rlabel metal2 48 1020 102 1073 0 Pixel_s1[0]
<< end >>
