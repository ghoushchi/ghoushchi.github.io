magic
tech scmos
timestamp 951572636
<< nwell >>
rect -6 53 42 105
rect 26 50 42 53
<< polysilicon >>
rect 11 97 13 99
rect 19 97 21 99
rect 27 97 29 99
rect 35 97 37 99
rect 11 80 13 89
rect 19 80 21 89
rect 2 78 21 80
rect 2 75 4 78
rect 0 55 2 75
rect 11 70 13 72
rect 19 70 21 72
rect -3 53 2 55
rect 27 56 29 57
rect 27 54 31 56
rect -3 45 -1 53
rect 11 51 13 54
rect 19 51 21 54
rect 29 52 31 54
rect 35 52 37 57
rect 9 49 13 51
rect 9 47 14 49
rect 18 47 22 51
rect 29 50 37 52
rect -3 43 2 45
rect 0 40 2 43
rect 12 44 14 47
rect 12 42 17 44
rect 0 38 13 40
rect 11 32 13 38
rect 15 32 17 42
rect 19 32 21 47
rect 29 44 31 50
rect 29 31 31 40
rect 27 29 37 31
rect 27 28 29 29
rect 35 28 37 29
rect 11 6 13 8
rect 15 6 17 8
rect 19 6 21 8
rect 27 6 29 8
rect 35 6 37 8
<< ndiffusion >>
rect 10 8 11 32
rect 13 8 15 32
rect 17 8 19 32
rect 21 8 22 32
rect 26 8 27 28
rect 29 8 30 28
rect 34 8 35 28
rect 37 8 38 28
<< pdiffusion >>
rect 10 89 11 97
rect 13 89 14 97
rect 18 89 19 97
rect 21 89 22 97
rect 10 54 11 70
rect 13 54 14 70
rect 18 54 19 70
rect 21 54 22 70
rect 26 57 27 97
rect 29 57 30 97
rect 34 57 35 97
rect 37 57 38 97
<< metal1 >>
rect -1 79 2 106
rect 5 103 13 105
rect 10 101 13 103
rect 6 97 10 99
rect 22 97 26 99
rect 38 97 42 99
rect 6 70 10 89
rect 14 70 18 89
rect 4 47 5 51
rect 13 47 17 54
rect 22 51 26 54
rect 30 53 34 57
rect 30 50 38 53
rect 14 44 18 47
rect 5 40 27 44
rect 5 33 9 40
rect 34 35 38 50
rect 6 32 10 33
rect -6 6 -2 8
rect 22 6 26 8
rect 30 31 38 35
rect 30 28 34 31
rect 30 1 33 8
rect 38 6 42 8
rect 29 -2 33 1
<< metal2 >>
rect 13 103 17 105
rect -6 99 5 103
rect 10 99 22 103
rect 26 99 38 103
rect -6 47 0 51
rect 4 47 42 51
rect -2 2 22 6
rect 26 2 38 6
<< ntransistor >>
rect 11 8 13 32
rect 15 8 17 32
rect 19 8 21 32
rect 27 8 29 28
rect 35 8 37 28
<< ptransistor >>
rect 11 89 13 97
rect 19 89 21 97
rect 11 54 13 70
rect 19 54 21 70
rect 27 57 29 97
rect 35 57 37 97
<< polycontact >>
rect -2 75 2 79
rect 5 47 9 51
rect 22 47 26 51
rect 27 40 31 44
<< ndcontact >>
rect 6 8 10 32
rect 22 8 26 32
rect 30 8 34 28
rect 38 8 42 28
<< pdcontact >>
rect 6 89 10 97
rect 14 89 18 97
rect 6 54 10 70
rect 14 54 18 70
rect 22 54 26 97
rect 30 57 34 97
rect 38 57 42 97
<< m2contact >>
rect 5 99 10 103
rect 22 99 26 103
rect 38 99 42 103
rect 0 47 4 51
rect -6 2 -2 6
rect 22 2 26 6
rect 38 2 42 6
<< psubstratepcontact >>
rect -6 8 -2 37
<< nsubstratencontact >>
rect 13 101 17 105
<< labels >>
rlabel metal1 0 99 0 99 1 clock
rlabel metal2 -5 49 -5 49 7 qual
rlabel metal2 6 3 6 3 4 Gnd
rlabel metal1 31 -1 31 -1 1 wordline
rlabel metal2 32 101 32 101 2 Vdd
<< end >>
