magic
tech scmos
timestamp 951381780
<< nwell >>
rect 615 1022 703 1056
<< polysilicon >>
rect 629 1046 631 1048
rect 637 1046 639 1048
rect 661 1046 663 1048
rect 669 1046 671 1048
rect 677 1046 679 1048
rect 685 1046 687 1048
rect 621 1036 623 1045
rect 653 1036 655 1045
rect 693 1036 695 1045
rect 621 1024 623 1026
rect 620 1022 623 1024
rect 629 1025 631 1026
rect 637 1025 639 1026
rect 629 1023 639 1025
rect 620 1012 622 1022
rect 629 1012 631 1023
rect 653 1013 655 1026
rect 661 1025 663 1026
rect 669 1025 671 1026
rect 661 1023 671 1025
rect 677 1025 679 1026
rect 685 1025 687 1026
rect 677 1023 687 1025
rect 661 1020 663 1023
rect 662 1016 663 1020
rect 685 1020 687 1023
rect 685 1016 686 1020
rect 661 1014 671 1016
rect 661 1013 663 1014
rect 669 1013 671 1014
rect 677 1014 687 1016
rect 677 1013 679 1014
rect 685 1013 687 1014
rect 693 1013 695 1026
rect 620 1010 623 1012
rect 621 1009 623 1010
rect 629 1010 639 1012
rect 629 1009 631 1010
rect 637 1009 639 1010
rect 621 1002 623 1004
rect 653 1006 655 1008
rect 693 1006 695 1008
rect 661 1001 663 1003
rect 669 1001 671 1003
rect 677 1001 679 1003
rect 685 1001 687 1003
rect 629 997 631 999
rect 637 997 639 999
<< ndiffusion >>
rect 620 1004 621 1009
rect 623 1004 624 1009
rect 628 999 629 1009
rect 631 999 632 1009
rect 636 999 637 1009
rect 639 999 640 1009
rect 652 1008 653 1013
rect 655 1008 656 1013
rect 660 1003 661 1013
rect 663 1003 664 1013
rect 668 1003 669 1013
rect 671 1003 672 1013
rect 676 1003 677 1013
rect 679 1003 680 1013
rect 684 1003 685 1013
rect 687 1003 688 1013
rect 692 1008 693 1013
rect 695 1008 696 1013
<< pdiffusion >>
rect 620 1026 621 1036
rect 623 1026 624 1036
rect 628 1026 629 1046
rect 631 1026 632 1046
rect 636 1026 637 1046
rect 639 1026 640 1046
rect 652 1026 653 1036
rect 655 1026 656 1036
rect 660 1026 661 1046
rect 663 1026 664 1046
rect 668 1026 669 1046
rect 671 1026 672 1046
rect 676 1026 677 1046
rect 679 1026 680 1046
rect 684 1026 685 1046
rect 687 1026 688 1046
rect 692 1026 693 1036
rect 695 1026 696 1036
<< metal1 >>
rect 617 1045 621 1056
rect 624 1046 628 1049
rect 640 1046 644 1049
rect 649 1045 653 1056
rect 656 1053 661 1056
rect 660 1052 661 1053
rect 671 1053 676 1056
rect 671 1052 672 1053
rect 656 1046 660 1049
rect 672 1046 676 1049
rect 688 1046 692 1049
rect 695 1045 699 1056
rect 616 1019 620 1026
rect 616 1015 625 1019
rect 616 1009 620 1015
rect 632 1009 636 1026
rect 648 1020 652 1026
rect 624 995 628 999
rect 620 991 624 995
rect 632 990 636 999
rect 640 1009 644 1014
rect 648 1016 658 1020
rect 648 1013 652 1016
rect 665 1013 668 1026
rect 656 1002 660 1003
rect 644 999 660 1002
rect 640 998 660 999
rect 672 1013 676 1014
rect 680 1013 683 1026
rect 696 1020 700 1026
rect 690 1016 700 1020
rect 696 1013 700 1016
rect 664 1000 668 1003
rect 680 1000 684 1003
rect 640 995 644 998
rect 664 997 672 1000
rect 668 990 672 997
rect 675 997 684 1000
rect 675 990 679 997
rect 688 995 692 1003
<< metal2 >>
rect 615 1053 703 1056
rect 615 1049 624 1053
rect 628 1049 640 1053
rect 644 1049 656 1053
rect 660 1049 672 1053
rect 676 1049 688 1053
rect 692 1049 703 1053
rect 644 1014 672 1018
rect 615 991 624 995
rect 628 991 640 995
rect 644 991 688 995
rect 692 991 703 995
rect 615 990 703 991
<< ntransistor >>
rect 621 1004 623 1009
rect 629 999 631 1009
rect 637 999 639 1009
rect 653 1008 655 1013
rect 661 1003 663 1013
rect 669 1003 671 1013
rect 677 1003 679 1013
rect 685 1003 687 1013
rect 693 1008 695 1013
<< ptransistor >>
rect 621 1026 623 1036
rect 629 1026 631 1046
rect 637 1026 639 1046
rect 653 1026 655 1036
rect 661 1026 663 1046
rect 669 1026 671 1046
rect 677 1026 679 1046
rect 685 1026 687 1046
rect 693 1026 695 1036
<< polycontact >>
rect 617 1041 621 1045
rect 649 1041 653 1045
rect 695 1041 699 1045
rect 625 1015 629 1019
rect 658 1016 662 1020
rect 686 1016 690 1020
<< ndcontact >>
rect 616 1004 620 1009
rect 624 999 628 1009
rect 632 999 636 1009
rect 640 999 644 1009
rect 648 1008 652 1013
rect 656 1003 660 1013
rect 664 1003 668 1013
rect 672 1003 676 1013
rect 680 1003 684 1013
rect 688 1003 692 1013
rect 696 1008 700 1013
<< pdcontact >>
rect 616 1026 620 1036
rect 624 1026 628 1046
rect 632 1026 636 1046
rect 640 1026 644 1046
rect 648 1026 652 1036
rect 656 1026 660 1046
rect 664 1026 668 1046
rect 672 1026 676 1046
rect 680 1026 684 1046
rect 688 1026 692 1046
rect 696 1026 700 1036
<< m2contact >>
rect 624 1049 628 1053
rect 640 1049 644 1053
rect 656 1049 660 1053
rect 672 1049 676 1053
rect 688 1049 692 1053
rect 624 991 628 995
rect 640 1014 644 1018
rect 672 1014 676 1018
rect 640 991 644 995
rect 688 991 692 995
<< psubstratepcontact >>
rect 616 991 620 1000
<< nsubstratencontact >>
rect 661 1052 671 1056
<< labels >>
rlabel metal2 634 1051 634 1051 1 Vdd
rlabel metal1 619 1052 619 1052 1 cntrl0
rlabel metal2 646 994 646 994 2 Gnd
rlabel metal1 651 1053 651 1053 1 cntrl1
rlabel metal1 697 1053 697 1053 1 cntrl2
rlabel metal1 669 997 669 997 2 buff1
rlabel metal1 676 997 676 997 2 buff2
rlabel metal1 633 997 633 997 3 buff0
<< end >>
