magic
tech scmos
timestamp 951112323
<< metal1 >>
rect 8 64 11 72
rect 15 64 18 68
rect 116 64 119 72
rect 123 64 126 68
rect 60 -373 64 -369
<< metal2 >>
rect 48 112 117 117
rect 152 112 164 117
rect 7 80 11 84
rect 115 80 119 84
rect 31 59 37 64
rect 0 25 5 29
rect 1 -25 5 -21
rect 1 -145 5 -141
rect 1 -335 4 -331
rect 28 -361 35 -355
rect 1 -385 6 -381
rect 1 -420 5 -415
<< m2contact >>
rect 8 72 12 76
rect 116 72 120 76
use inverters inverters_0
timestamp 951078626
transform 1 0 46 0 1 72
box -37 -12 2 45
use inverters inverters_1
timestamp 951078626
transform 1 0 154 0 1 72
box -37 -12 2 45
use SetCell SetCell_0
timestamp 951088720
transform 1 0 17 0 1 3
box -17 -3 147 61
use ResetCell ResetCell_0
timestamp 951088720
transform 1 0 22 0 -1 -9
box -21 -13 142 51
use ResetCellflip ResetCellflip_0
timestamp 951112323
transform 1 0 -8 0 1 -207
box 9 87 172 151
use ResetCell ResetCell_1
timestamp 951088720
transform 1 0 22 0 -1 -129
box -21 -13 142 51
use ResetCellflip ResetCellflip_1
timestamp 951112323
transform 1 0 -8 0 1 -327
box 9 87 172 151
use ResetCell ResetCell_2
timestamp 951088720
transform 1 0 22 0 -1 -249
box -21 -13 142 51
use ResetCellflip ResetCellflip_2
timestamp 951112323
transform 1 0 -8 0 1 -447
box 9 87 172 151
use ResetCell ResetCell_3
timestamp 951088720
transform 1 0 22 0 -1 -369
box -21 -13 142 51
<< labels >>
rlabel metal2 34 62 34 62 5 Vdd
rlabel metal2 31 -358 31 -358 1 Gnd
rlabel metal2 2 -384 2 -384 3 Pix_Mux_s1[0]
rlabel metal2 2 -334 2 -334 3 Pix_Mux_s1[1]
rlabel space 2 -264 2 -264 3 Pix_Mux_s1[2]
rlabel space 2 -214 2 -214 3 Pix_Mux_s1[3]
rlabel metal2 2 -144 2 -144 3 Pix_Mux_s1[4]
rlabel space 2 -94 2 -94 3 Pix_Mux_s1[5]
rlabel metal2 2 -24 2 -24 3 Pix_Mux_s1[6]
rlabel metal2 1 26 1 26 3 Pix_Mux_s1[7]
rlabel metal2 8 82 8 82 1 Phi2
rlabel metal2 116 82 116 82 1 c8_Phi1_q1
<< end >>
