magic
tech scmos
timestamp 951219335
<< error_p >>
rect 4 40 5 41
rect -1 35 0 40
rect 4 38 15 40
rect 4 34 5 35
rect 14 34 15 38
rect 17 35 18 40
rect 4 19 5 22
<< pwell >>
rect 0 0 32 29
<< nwell >>
rect 0 29 32 45
<< polysilicon >>
rect 5 38 9 40
rect 23 38 27 40
rect 5 33 9 35
rect 5 22 7 33
rect 23 32 27 35
rect 12 30 27 32
rect 5 21 18 22
rect 5 20 20 21
rect 5 19 7 20
rect 25 19 27 30
rect 5 9 7 11
rect 15 7 19 8
rect 25 9 27 11
rect 0 5 8 7
rect 12 5 20 7
rect 24 5 32 7
<< ndiffusion >>
rect 0 19 4 22
rect 28 19 32 22
rect 4 15 5 19
rect 0 11 5 15
rect 7 15 8 19
rect 7 11 12 15
rect 24 15 25 19
rect 8 7 12 11
rect 20 11 25 15
rect 27 15 28 19
rect 27 11 32 15
rect 20 7 24 11
rect 8 4 12 5
rect 20 4 24 5
<< pdiffusion >>
rect 0 38 4 41
rect 28 38 32 41
rect 4 35 5 38
rect 9 35 10 38
rect 22 35 23 38
rect 27 35 28 38
<< metal1 >>
rect 4 41 28 45
rect 0 38 4 41
rect 28 38 32 41
rect 10 32 14 34
rect 0 26 4 27
rect 0 19 4 22
rect 8 30 14 32
rect 8 26 10 30
rect 8 19 12 26
rect 18 25 22 34
rect 28 26 32 27
rect 22 21 24 25
rect 20 19 24 21
rect 28 19 32 22
rect 0 9 15 12
rect 19 9 32 12
rect 7 0 8 4
rect 19 0 20 4
<< metal2 >>
rect 0 31 4 45
rect 10 30 13 45
rect 0 8 4 27
rect 8 27 13 30
rect 8 4 11 27
rect 19 20 22 45
rect 16 17 22 20
rect 28 31 32 45
rect 16 4 19 17
rect 28 12 32 27
rect 7 0 11 4
rect 23 8 32 12
rect 23 0 27 8
<< ntransistor >>
rect 5 11 7 19
rect 25 11 27 19
rect 8 5 12 7
rect 20 5 24 7
<< ptransistor >>
rect 5 35 9 38
rect 23 35 27 38
<< polycontact >>
rect 10 26 14 30
rect 18 21 22 25
rect 15 8 19 12
<< ndcontact >>
rect 0 15 4 19
rect 8 15 12 19
rect 20 15 24 19
rect 28 15 32 19
rect 8 0 12 4
rect 20 0 24 4
<< pdcontact >>
rect 0 34 4 38
rect 10 34 14 38
rect 18 34 22 38
rect 28 34 32 38
<< m2contact >>
rect 0 27 4 31
rect 28 27 32 31
rect 3 0 7 4
rect 15 0 19 4
<< psubstratepcontact >>
rect 0 22 4 26
rect 28 22 32 26
<< nsubstratencontact >>
rect 0 41 4 45
rect 28 41 32 45
<< labels >>
rlabel metal1 22 43 22 43 1 Vdd
rlabel metal2 20 40 20 40 1 bit_b
rlabel metal2 12 40 12 40 1 bit
rlabel m2contact 30 29 30 29 1 gnd
rlabel metal1 9 31 9 31 1 a
rlabel m2contact 2 29 2 29 1 gnda
rlabel metal1 20 30 20 30 5 a_b
<< end >>
