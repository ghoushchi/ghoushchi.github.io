magic
tech scmos
timestamp 951727448
<< pwell >>
rect 0 0 56 32
<< nwell >>
rect 0 32 56 64
<< polysilicon >>
rect 15 60 45 62
rect 11 56 13 58
rect 15 56 17 60
rect 23 56 25 58
rect 27 56 29 58
rect 43 52 45 60
rect 43 46 45 48
rect 43 44 46 46
rect 11 23 13 40
rect 15 38 17 40
rect 23 37 25 40
rect 27 39 29 40
rect 27 37 37 39
rect 19 33 20 36
rect 24 35 25 37
rect 19 23 21 33
rect 35 29 37 37
rect 44 34 46 44
rect 27 27 37 29
rect 43 32 46 34
rect 27 23 29 27
rect 35 23 37 25
rect 11 9 13 11
rect 19 9 21 11
rect 27 9 29 11
rect 35 9 37 11
rect 43 9 45 32
rect 35 7 45 9
<< ndiffusion >>
rect 10 11 11 23
rect 13 11 14 23
rect 18 11 19 23
rect 21 22 27 23
rect 21 18 22 22
rect 26 18 27 22
rect 21 11 27 18
rect 29 11 30 23
rect 34 11 35 23
rect 37 11 38 23
<< pdiffusion >>
rect 10 40 11 56
rect 13 40 15 56
rect 17 53 23 56
rect 17 41 18 53
rect 22 41 23 53
rect 17 40 23 41
rect 25 40 27 56
rect 29 40 30 56
<< metal1 >>
rect 0 58 46 60
rect 0 56 34 58
rect 14 41 18 49
rect 7 30 10 31
rect 14 30 17 41
rect 38 56 46 58
rect 50 56 56 60
rect 45 48 46 52
rect 38 36 41 37
rect 24 33 30 36
rect 14 27 22 30
rect 22 22 26 26
rect 46 25 50 27
rect 22 17 26 18
rect 18 11 30 14
rect 6 8 10 11
rect 38 8 42 11
rect 0 5 46 8
rect 50 5 56 8
rect 0 4 56 5
<< ntransistor >>
rect 11 11 13 23
rect 19 11 21 23
rect 27 11 29 23
rect 35 11 37 23
<< ptransistor >>
rect 11 40 13 56
rect 15 40 17 56
rect 23 40 25 56
rect 27 40 29 56
<< polycontact >>
rect 41 48 45 52
rect 7 31 11 35
rect 37 37 41 41
rect 20 33 24 37
<< ndcontact >>
rect 6 11 10 23
rect 14 11 18 23
rect 22 18 26 22
rect 30 11 34 23
rect 38 11 42 23
<< pdcontact >>
rect 6 40 10 56
rect 18 41 22 53
rect 30 40 34 56
<< m2contact >>
rect 6 26 10 30
rect 46 48 50 52
rect 30 32 34 36
rect 38 32 42 36
rect 22 26 26 30
<< psubstratepcontact >>
rect 46 5 50 25
<< nsubstratencontact >>
rect 34 46 38 58
rect 46 56 50 60
<< psubstratepdiff >>
rect 46 25 50 27
rect 46 4 50 5
<< labels >>
rlabel m2contact 8 28 8 28 6 In2
rlabel m2contact 24 28 24 28 6 Out_b
rlabel m2contact 32 34 32 34 6 In0
rlabel m2contact 40 34 40 34 6 In1
rlabel metal1 52 58 52 58 6 Vdd
rlabel metal1 4 58 4 58 6 Vdd
rlabel metal1 52 6 52 6 6 GND
rlabel metal1 4 6 4 6 6 GND
rlabel m2contact 48 50 48 50 6 In3
<< end >>
