magic
tech scmos
timestamp 950486748
<< polysilicon >>
rect 165 127 167 129
rect 175 127 177 129
rect 183 127 185 129
rect 193 127 195 129
rect 201 127 203 129
rect 211 127 213 129
rect 219 127 221 129
rect 229 127 231 129
rect 237 127 239 129
rect 247 127 249 129
rect 165 112 167 113
rect 166 110 167 112
rect 175 110 177 111
rect 183 110 185 111
rect 193 110 195 111
rect 201 110 203 111
rect 211 110 213 111
rect 219 110 221 111
rect 229 110 231 111
rect 237 110 239 111
rect 247 110 249 111
rect 166 108 249 110
rect 12 96 14 98
rect 20 97 30 99
rect 20 96 22 97
rect 28 96 30 97
rect 36 96 38 98
rect 52 94 54 96
rect 60 94 62 97
rect 12 85 14 86
rect 20 85 22 86
rect 12 83 22 85
rect 28 85 30 86
rect 36 85 38 86
rect 28 83 38 85
rect 52 83 54 84
rect 60 83 62 84
rect 52 81 62 83
rect 112 96 114 98
rect 120 97 130 99
rect 120 96 122 97
rect 128 96 130 97
rect 136 96 138 99
rect 156 96 158 98
rect 164 96 166 98
rect 172 96 174 98
rect 85 93 87 95
rect 98 93 101 95
rect 99 92 101 93
rect 99 89 100 92
rect 120 84 122 86
rect 128 85 130 86
rect 112 83 114 84
rect 128 83 132 85
rect 108 81 114 83
rect 136 83 138 86
rect 156 83 158 84
rect 164 83 166 84
rect 172 83 174 84
rect 156 81 182 83
rect 87 66 108 67
rect 91 62 104 66
rect 136 64 165 68
rect 87 61 108 62
rect 12 46 14 48
rect 20 46 22 48
rect 28 46 30 48
rect 36 46 38 49
rect 52 47 62 49
rect 85 49 94 51
rect 85 48 87 49
rect 52 46 54 47
rect 60 46 62 47
rect 12 21 14 22
rect 20 21 22 22
rect 28 21 30 22
rect 36 21 38 22
rect 12 19 38 21
rect 52 20 54 22
rect 60 20 62 22
rect 106 46 108 49
rect 112 47 124 49
rect 114 46 116 47
rect 122 46 124 47
rect 142 47 154 49
rect 166 49 179 51
rect 142 46 144 47
rect 150 46 152 47
rect 158 46 160 49
rect 166 48 168 49
rect 193 49 267 51
rect 193 48 195 49
rect 201 48 203 49
rect 209 48 211 49
rect 217 48 219 49
rect 225 48 227 49
rect 233 48 235 49
rect 241 48 243 49
rect 249 48 251 49
rect 257 48 259 49
rect 265 48 267 49
rect 85 22 87 24
rect 106 22 108 24
rect 114 22 116 24
rect 122 22 124 24
rect 142 22 144 24
rect 150 22 152 24
rect 158 22 160 24
rect 166 22 168 24
rect 193 22 195 24
rect 201 22 203 24
rect 209 22 211 24
rect 217 22 219 24
rect 225 22 227 24
rect 233 22 235 24
rect 241 22 243 24
rect 249 22 251 24
rect 257 22 259 24
rect 265 22 267 24
<< ndiffusion >>
rect 0 314 8 315
rect 0 142 1 314
rect 5 307 8 314
rect 32 307 34 315
rect 5 289 6 307
rect 9 302 30 303
rect 9 294 11 302
rect 27 294 30 302
rect 9 293 30 294
rect 9 292 20 293
rect 5 288 16 289
rect 5 280 7 288
rect 15 280 16 288
rect 5 279 16 280
rect 5 265 6 279
rect 19 277 20 292
rect 28 277 30 293
rect 19 276 30 277
rect 9 274 30 276
rect 9 270 11 274
rect 27 270 30 274
rect 9 269 30 270
rect 9 268 20 269
rect 5 263 16 265
rect 5 259 6 263
rect 14 259 16 263
rect 5 258 16 259
rect 5 246 6 258
rect 19 255 20 268
rect 9 254 20 255
rect 9 250 11 254
rect 19 250 20 254
rect 9 249 20 250
rect 5 245 16 246
rect 5 241 7 245
rect 15 241 16 245
rect 5 240 16 241
rect 5 222 6 240
rect 19 237 20 249
rect 28 237 30 269
rect 9 235 30 237
rect 9 227 11 235
rect 27 227 30 235
rect 9 225 30 227
rect 5 221 16 222
rect 5 213 7 221
rect 15 213 16 221
rect 5 212 16 213
rect 5 198 6 212
rect 19 209 20 225
rect 28 209 30 225
rect 9 207 30 209
rect 9 203 11 207
rect 27 203 30 207
rect 9 201 30 203
rect 19 200 30 201
rect 5 197 16 198
rect 5 193 7 197
rect 15 193 16 197
rect 5 192 16 193
rect 5 174 6 192
rect 19 189 20 200
rect 9 188 20 189
rect 28 188 30 200
rect 9 187 30 188
rect 9 179 11 187
rect 27 179 30 187
rect 9 177 30 179
rect 5 173 16 174
rect 5 165 7 173
rect 15 165 16 173
rect 5 164 16 165
rect 19 161 20 177
rect 9 160 20 161
rect 9 156 10 160
rect 18 157 20 160
rect 28 157 30 177
rect 18 156 30 157
rect 9 155 30 156
rect 9 151 10 155
rect 18 151 20 155
rect 28 151 30 155
rect 9 150 30 151
rect 33 203 34 307
rect 42 203 43 315
rect 33 171 43 203
rect 33 147 34 171
rect 5 146 34 147
rect 5 142 6 146
rect 14 143 34 146
rect 42 143 43 171
rect 14 142 43 143
rect 0 141 43 142
rect 242 203 243 315
rect 251 307 254 315
rect 278 314 285 315
rect 278 307 280 314
rect 251 203 252 307
rect 242 170 252 203
rect 242 142 243 170
rect 251 147 252 170
rect 255 302 276 303
rect 255 294 258 302
rect 274 294 276 302
rect 255 293 276 294
rect 255 277 257 293
rect 265 292 276 293
rect 265 277 266 292
rect 279 289 280 307
rect 269 288 280 289
rect 269 280 270 288
rect 278 280 280 288
rect 269 279 280 280
rect 255 276 266 277
rect 255 274 276 276
rect 255 270 258 274
rect 274 270 276 274
rect 255 268 276 270
rect 255 236 257 268
rect 265 255 266 268
rect 279 265 280 279
rect 269 263 280 265
rect 269 259 271 263
rect 279 259 280 263
rect 269 258 280 259
rect 265 254 276 255
rect 265 250 266 254
rect 274 250 276 254
rect 265 249 276 250
rect 265 237 266 249
rect 279 246 280 258
rect 269 245 280 246
rect 269 241 270 245
rect 278 241 280 245
rect 269 240 280 241
rect 265 236 276 237
rect 255 235 276 236
rect 255 227 258 235
rect 274 227 276 235
rect 255 225 276 227
rect 255 209 257 225
rect 265 209 266 225
rect 279 222 280 240
rect 269 221 280 222
rect 269 213 270 221
rect 278 213 280 221
rect 269 212 280 213
rect 255 207 276 209
rect 255 203 258 207
rect 274 203 276 207
rect 255 201 276 203
rect 255 200 266 201
rect 255 188 257 200
rect 265 189 266 200
rect 279 198 280 212
rect 269 197 280 198
rect 269 193 270 197
rect 278 193 280 197
rect 269 192 280 193
rect 265 188 276 189
rect 255 187 276 188
rect 255 179 258 187
rect 274 179 276 187
rect 255 177 276 179
rect 255 165 257 177
rect 265 165 266 177
rect 279 174 280 192
rect 255 164 266 165
rect 269 173 280 174
rect 269 165 270 173
rect 278 165 280 173
rect 269 164 280 165
rect 255 156 257 164
rect 265 161 266 164
rect 265 160 276 161
rect 265 156 267 160
rect 275 156 276 160
rect 255 155 276 156
rect 255 151 257 155
rect 265 151 267 155
rect 275 151 276 155
rect 255 150 276 151
rect 279 154 280 164
rect 284 154 285 314
rect 279 147 285 154
rect 251 146 285 147
rect 251 142 252 146
rect 256 142 275 146
rect 283 142 285 146
rect 242 141 285 142
rect 28 109 111 129
rect 164 116 165 127
rect 160 113 165 116
rect 167 124 175 127
rect 167 113 169 124
rect 168 112 169 113
rect 173 112 175 124
rect 168 111 175 112
rect 177 124 183 127
rect 177 112 178 124
rect 182 112 183 124
rect 177 111 183 112
rect 185 124 193 127
rect 185 112 187 124
rect 191 112 193 124
rect 185 111 193 112
rect 195 124 201 127
rect 195 112 196 124
rect 200 112 201 124
rect 195 111 201 112
rect 203 124 211 127
rect 203 112 205 124
rect 209 112 211 124
rect 203 111 211 112
rect 213 124 219 127
rect 213 112 214 124
rect 218 112 219 124
rect 213 111 219 112
rect 221 124 229 127
rect 221 112 223 124
rect 227 112 229 124
rect 221 111 229 112
rect 231 124 237 127
rect 231 112 232 124
rect 236 112 237 124
rect 231 111 237 112
rect 239 124 247 127
rect 239 112 241 124
rect 245 112 247 124
rect 239 111 247 112
rect 249 124 254 127
rect 249 112 250 124
rect 249 111 254 112
rect 11 88 12 96
rect 7 86 12 88
rect 14 88 15 96
rect 19 88 20 96
rect 14 86 20 88
rect 22 88 23 96
rect 27 88 28 96
rect 22 86 28 88
rect 30 88 31 96
rect 35 88 36 96
rect 30 86 36 88
rect 38 88 39 96
rect 38 86 43 88
rect 51 87 52 94
rect 47 84 52 87
rect 54 92 60 94
rect 54 84 55 92
rect 59 84 60 92
rect 62 92 67 94
rect 62 84 63 92
rect 87 95 98 96
rect 87 92 98 93
rect 95 90 98 92
rect 111 88 112 96
rect 109 84 112 88
rect 114 84 115 96
rect 119 86 120 96
rect 122 90 128 96
rect 122 86 123 90
rect 127 86 128 90
rect 130 88 131 96
rect 135 88 136 96
rect 130 86 136 88
rect 138 90 143 96
rect 138 86 139 90
rect 155 84 156 96
rect 158 90 164 96
rect 158 86 159 90
rect 163 86 164 90
rect 158 84 164 86
rect 166 92 167 96
rect 171 92 172 96
rect 166 84 172 92
rect 174 84 175 96
<< pdiffusion >>
rect 214 80 271 81
rect 222 64 255 80
rect 214 63 271 64
rect 11 22 12 46
rect 14 22 15 46
rect 19 22 20 46
rect 22 22 23 46
rect 27 22 28 46
rect 30 22 31 46
rect 35 22 36 46
rect 38 40 43 46
rect 38 22 39 40
rect 51 22 52 46
rect 54 22 55 46
rect 59 22 60 46
rect 62 42 67 46
rect 62 22 63 42
rect 84 24 85 48
rect 87 44 90 48
rect 161 46 166 48
rect 101 45 106 46
rect 87 24 88 44
rect 105 25 106 45
rect 101 24 106 25
rect 108 36 114 46
rect 108 24 109 36
rect 113 24 114 36
rect 116 44 122 46
rect 116 32 117 44
rect 121 32 122 44
rect 116 24 122 32
rect 124 45 129 46
rect 124 25 125 45
rect 124 24 129 25
rect 141 30 142 46
rect 137 24 142 30
rect 144 36 150 46
rect 144 24 145 36
rect 149 24 150 36
rect 152 44 158 46
rect 152 32 153 44
rect 157 32 158 44
rect 152 24 158 32
rect 160 45 166 46
rect 160 25 161 45
rect 165 25 166 45
rect 160 24 166 25
rect 168 43 171 48
rect 188 44 193 48
rect 168 41 178 43
rect 168 25 174 41
rect 168 24 178 25
rect 192 24 193 44
rect 195 28 196 48
rect 200 28 201 48
rect 195 24 201 28
rect 203 24 204 48
rect 208 24 209 48
rect 211 28 212 48
rect 216 28 217 48
rect 211 24 217 28
rect 219 24 220 48
rect 224 24 225 48
rect 227 28 228 48
rect 232 28 233 48
rect 227 24 233 28
rect 235 24 236 48
rect 240 24 241 48
rect 243 28 244 48
rect 248 28 249 48
rect 243 24 249 28
rect 251 24 252 48
rect 256 24 257 48
rect 259 28 260 48
rect 264 28 265 48
rect 259 24 265 28
rect 267 24 268 48
<< metal1 >>
rect 0 314 8 315
rect 0 142 1 314
rect 5 307 8 314
rect 32 307 34 315
rect 5 289 6 307
rect 10 302 29 303
rect 10 294 11 302
rect 27 294 29 302
rect 10 293 29 294
rect 5 288 16 289
rect 5 280 7 288
rect 15 280 16 288
rect 5 279 16 280
rect 5 264 6 279
rect 28 277 29 293
rect 20 275 29 277
rect 10 274 29 275
rect 10 270 11 274
rect 27 270 29 274
rect 10 269 29 270
rect 5 263 15 264
rect 5 259 6 263
rect 14 259 15 263
rect 5 258 15 259
rect 5 246 6 258
rect 10 254 20 255
rect 10 250 11 254
rect 19 250 20 254
rect 10 249 20 250
rect 5 245 16 246
rect 5 241 7 245
rect 15 241 16 245
rect 5 240 16 241
rect 5 222 6 240
rect 28 237 29 269
rect 20 236 29 237
rect 10 235 29 236
rect 10 227 11 235
rect 27 227 29 235
rect 10 226 29 227
rect 20 225 29 226
rect 5 221 16 222
rect 5 213 7 221
rect 15 213 16 221
rect 5 212 16 213
rect 5 198 6 212
rect 28 209 29 225
rect 20 208 29 209
rect 10 207 29 208
rect 10 203 11 207
rect 27 203 29 207
rect 33 203 34 307
rect 42 203 43 315
rect 10 202 29 203
rect 20 200 29 202
rect 5 197 16 198
rect 5 193 7 197
rect 15 193 16 197
rect 5 192 16 193
rect 5 174 6 192
rect 28 198 29 200
rect 67 198 219 320
rect 242 203 243 315
rect 251 307 254 315
rect 278 314 285 315
rect 278 307 280 314
rect 251 203 252 307
rect 256 302 275 303
rect 256 294 258 302
rect 274 294 275 302
rect 256 293 275 294
rect 256 277 257 293
rect 279 289 280 307
rect 269 288 280 289
rect 269 280 270 288
rect 278 280 280 288
rect 269 279 280 280
rect 256 275 265 277
rect 256 274 275 275
rect 256 270 258 274
rect 274 270 275 274
rect 256 269 275 270
rect 256 268 265 269
rect 256 236 257 268
rect 279 264 280 279
rect 270 263 280 264
rect 270 259 271 263
rect 279 259 280 263
rect 270 258 280 259
rect 265 254 275 255
rect 265 250 266 254
rect 274 250 275 254
rect 265 249 275 250
rect 279 246 280 258
rect 269 245 280 246
rect 269 241 270 245
rect 278 241 280 245
rect 269 240 280 241
rect 256 235 275 236
rect 256 227 258 235
rect 274 227 275 235
rect 256 226 275 227
rect 256 225 265 226
rect 256 209 257 225
rect 279 222 280 240
rect 269 221 280 222
rect 269 213 270 221
rect 278 213 280 221
rect 269 212 280 213
rect 256 208 265 209
rect 256 207 275 208
rect 256 203 258 207
rect 274 203 275 207
rect 256 202 275 203
rect 256 200 265 202
rect 256 198 257 200
rect 28 188 257 198
rect 279 198 280 212
rect 269 197 280 198
rect 269 193 270 197
rect 278 193 280 197
rect 269 192 280 193
rect 10 187 275 188
rect 10 179 11 187
rect 27 179 258 187
rect 274 179 275 187
rect 10 178 275 179
rect 20 177 265 178
rect 5 173 16 174
rect 5 165 7 173
rect 15 165 16 173
rect 18 157 20 160
rect 28 157 29 177
rect 18 156 29 157
rect 10 155 29 156
rect 18 151 20 155
rect 28 151 29 155
rect 5 146 15 147
rect 5 142 6 146
rect 14 142 15 146
rect 0 140 15 142
rect 0 104 2 140
rect 6 139 15 140
rect 6 104 7 139
rect 19 129 29 151
rect 33 171 43 172
rect 33 143 34 171
rect 42 143 43 171
rect 67 168 219 177
rect 242 170 252 172
rect 33 141 43 143
rect 242 142 243 170
rect 251 147 252 170
rect 256 165 257 177
rect 279 174 280 192
rect 256 164 265 165
rect 269 173 280 174
rect 269 165 270 173
rect 278 165 280 173
rect 269 164 280 165
rect 256 156 257 164
rect 265 160 276 161
rect 265 156 267 160
rect 275 156 276 160
rect 256 155 276 156
rect 256 151 257 155
rect 265 151 267 155
rect 279 154 280 164
rect 284 154 285 314
rect 251 146 257 147
rect 251 142 252 146
rect 256 142 257 146
rect 242 141 257 142
rect 33 139 254 141
rect 141 135 159 139
rect 163 136 178 139
rect 163 135 165 136
rect 182 136 196 139
rect 33 133 133 135
rect 137 131 138 135
rect 28 109 29 129
rect 70 109 111 112
rect 127 127 148 128
rect 152 127 153 131
rect 127 126 157 127
rect 127 122 148 126
rect 152 122 153 126
rect 127 118 157 122
rect 160 127 164 135
rect 169 132 174 133
rect 173 128 174 132
rect 169 124 174 128
rect 137 112 151 114
rect 173 112 174 124
rect 0 100 3 104
rect 27 100 29 104
rect 33 100 34 104
rect 42 100 43 104
rect 0 96 1 100
rect 5 96 10 100
rect 23 96 27 100
rect 0 95 7 96
rect 0 87 3 95
rect 7 87 11 88
rect 0 85 11 87
rect 0 81 1 85
rect 5 81 7 85
rect 11 81 12 85
rect 0 77 12 81
rect 8 75 12 77
rect 8 70 12 71
rect 16 62 19 88
rect 47 100 49 104
rect 53 100 55 104
rect 47 99 59 100
rect 47 96 55 99
rect 47 94 51 96
rect 70 98 73 109
rect 141 108 142 112
rect 146 108 147 112
rect 169 111 174 112
rect 178 124 182 135
rect 200 136 214 139
rect 137 105 158 108
rect 137 104 138 105
rect 77 100 78 104
rect 126 100 127 104
rect 66 95 73 98
rect 23 85 27 88
rect 23 80 27 81
rect 23 75 27 76
rect 23 70 27 71
rect 32 62 35 88
rect 46 87 47 88
rect 0 57 1 61
rect 5 57 8 61
rect 12 57 13 61
rect 0 56 13 57
rect 0 52 1 56
rect 5 52 7 56
rect 11 55 13 56
rect 16 59 35 62
rect 0 51 11 52
rect 0 47 7 51
rect 0 46 11 47
rect 16 46 19 59
rect 0 22 3 46
rect 23 51 27 52
rect 23 46 27 47
rect 32 46 35 59
rect 39 62 42 81
rect 46 80 50 87
rect 46 75 50 76
rect 46 70 50 71
rect 56 62 59 84
rect 62 80 66 84
rect 62 75 66 76
rect 62 70 66 71
rect 39 59 59 62
rect 39 51 42 59
rect 0 18 1 22
rect 5 18 10 22
rect 0 17 10 18
rect 23 17 27 22
rect 0 13 1 17
rect 5 13 6 17
rect 10 13 11 17
rect 47 46 51 52
rect 56 46 59 59
rect 70 51 73 95
rect 80 96 84 100
rect 102 99 111 100
rect 106 96 111 99
rect 162 96 165 108
rect 178 105 182 112
rect 186 132 192 133
rect 186 128 187 132
rect 191 128 192 132
rect 186 124 192 128
rect 186 112 187 124
rect 191 112 192 124
rect 186 111 192 112
rect 196 124 200 135
rect 218 136 232 139
rect 196 105 200 112
rect 204 132 210 133
rect 204 128 205 132
rect 209 128 210 132
rect 204 124 210 128
rect 204 112 205 124
rect 209 112 210 124
rect 204 111 210 112
rect 214 124 218 135
rect 236 136 250 139
rect 182 99 200 101
rect 106 95 107 96
rect 80 91 84 92
rect 80 86 84 87
rect 80 80 84 82
rect 80 74 84 76
rect 98 88 100 91
rect 87 66 90 88
rect 98 85 101 88
rect 94 82 101 85
rect 94 66 97 82
rect 105 66 108 81
rect 66 48 73 51
rect 78 56 82 57
rect 78 48 82 52
rect 39 40 41 44
rect 45 40 47 44
rect 0 12 10 13
rect 31 0 34 22
rect 39 20 43 22
rect 63 42 67 43
rect 39 17 46 20
rect 41 16 47 17
rect 41 13 42 16
rect 46 13 47 16
rect 55 0 58 22
rect 63 17 67 22
rect 65 13 67 17
rect 70 0 73 48
rect 88 44 91 62
rect 94 51 97 62
rect 105 52 108 62
rect 119 93 131 96
rect 135 93 151 96
rect 123 85 127 86
rect 143 86 144 90
rect 139 85 148 86
rect 105 51 111 52
rect 105 49 108 51
rect 80 20 84 24
rect 80 17 90 20
rect 80 13 81 17
rect 85 13 86 17
rect 80 12 90 13
rect 95 0 98 47
rect 115 46 118 84
rect 123 80 127 81
rect 123 74 127 76
rect 139 81 144 85
rect 155 93 167 96
rect 163 86 175 87
rect 159 84 175 86
rect 186 95 189 99
rect 193 97 200 99
rect 193 95 196 97
rect 196 92 200 93
rect 179 88 192 91
rect 132 68 135 81
rect 139 80 148 81
rect 143 76 144 80
rect 148 76 150 80
rect 139 75 148 76
rect 143 71 144 75
rect 159 68 162 84
rect 167 75 171 76
rect 179 78 185 81
rect 139 65 162 68
rect 139 60 142 65
rect 126 57 142 60
rect 179 66 182 78
rect 126 46 129 57
rect 133 46 137 50
rect 165 52 168 64
rect 101 45 105 46
rect 115 44 121 46
rect 115 42 117 44
rect 105 39 117 42
rect 101 24 105 25
rect 117 31 121 32
rect 125 45 129 46
rect 113 25 125 27
rect 136 42 137 46
rect 132 41 137 42
rect 136 37 137 41
rect 132 36 137 37
rect 136 32 137 36
rect 147 44 151 52
rect 155 51 171 52
rect 158 49 171 51
rect 161 45 165 46
rect 141 40 153 44
rect 129 25 145 27
rect 113 24 145 25
rect 149 25 161 27
rect 149 24 165 25
rect 168 0 171 49
rect 179 51 182 62
rect 189 53 192 88
rect 196 87 200 88
rect 196 82 200 83
rect 204 83 208 111
rect 214 105 218 112
rect 222 132 228 133
rect 222 128 223 132
rect 227 128 228 132
rect 222 124 228 128
rect 222 112 223 124
rect 227 112 228 124
rect 211 99 219 101
rect 211 95 213 99
rect 217 95 219 99
rect 211 94 219 95
rect 211 90 213 94
rect 217 90 219 94
rect 222 84 228 112
rect 232 124 236 135
rect 232 106 236 112
rect 232 99 236 102
rect 240 132 246 133
rect 240 128 241 132
rect 245 128 246 132
rect 240 124 246 128
rect 240 112 241 124
rect 245 112 246 124
rect 240 84 246 112
rect 250 124 254 135
rect 250 106 254 112
rect 250 99 254 102
rect 222 83 246 84
rect 204 80 249 83
rect 261 80 270 151
rect 279 147 285 154
rect 274 146 285 147
rect 274 142 275 146
rect 283 142 285 146
rect 274 140 285 142
rect 274 100 275 140
rect 279 137 285 140
rect 283 133 285 137
rect 279 132 285 133
rect 283 128 285 132
rect 279 127 285 128
rect 283 123 285 127
rect 279 122 285 123
rect 283 118 285 122
rect 279 117 285 118
rect 283 113 285 117
rect 279 112 285 113
rect 283 108 285 112
rect 279 107 285 108
rect 283 103 285 107
rect 279 100 285 103
rect 274 99 285 100
rect 278 95 279 99
rect 283 95 285 99
rect 204 78 214 80
rect 196 77 200 78
rect 211 65 214 78
rect 196 64 214 65
rect 222 73 249 80
rect 196 63 222 64
rect 196 61 217 63
rect 196 48 200 61
rect 174 41 179 43
rect 178 40 179 41
rect 183 40 184 44
rect 178 39 184 40
rect 178 35 179 39
rect 183 35 184 39
rect 178 34 184 35
rect 178 30 179 34
rect 183 30 184 34
rect 178 29 184 30
rect 178 25 179 29
rect 183 25 184 29
rect 174 24 184 25
rect 204 48 208 54
rect 211 48 217 61
rect 211 28 212 48
rect 216 28 217 48
rect 220 48 224 54
rect 227 48 233 73
rect 227 28 228 48
rect 232 28 233 48
rect 236 48 240 54
rect 243 55 249 73
rect 243 51 265 55
rect 243 48 249 51
rect 259 48 265 51
rect 243 28 244 48
rect 248 28 249 48
rect 259 28 260 48
rect 264 28 265 48
rect 268 51 272 54
rect 284 52 285 88
rect 276 51 285 52
rect 268 50 285 51
rect 268 49 276 50
rect 268 48 272 49
rect 175 20 179 24
rect 183 23 272 24
rect 183 20 188 23
rect 175 19 188 20
rect 192 19 196 23
rect 200 19 204 23
rect 208 19 212 23
rect 216 19 220 23
rect 224 19 228 23
rect 232 19 236 23
rect 240 19 244 23
rect 248 19 252 23
rect 256 19 260 23
rect 264 21 272 23
rect 276 45 280 46
rect 276 40 280 41
rect 276 35 280 36
rect 276 30 280 31
rect 276 25 280 26
rect 264 20 280 21
rect 264 19 276 20
rect 175 18 276 19
rect 178 14 184 18
rect 192 17 196 18
rect 200 17 204 18
rect 208 17 212 18
rect 216 17 220 18
rect 224 17 228 18
rect 232 17 236 18
rect 240 17 244 18
rect 248 17 252 18
rect 256 17 260 18
rect 264 17 268 18
rect 284 18 285 50
rect 280 16 285 18
rect 276 14 285 16
rect 271 12 285 14
<< metal2 >>
rect 68 315 218 319
rect 0 139 20 315
rect 68 173 72 315
rect 214 173 218 315
rect 68 169 218 173
rect 265 141 285 315
rect 0 136 11 139
rect 0 132 2 136
rect 6 135 11 136
rect 15 135 20 139
rect 262 137 285 141
rect 6 132 20 135
rect 0 128 20 132
rect 0 124 2 128
rect 6 124 20 128
rect 0 116 20 124
rect 132 131 133 135
rect 137 131 138 135
rect 142 131 144 135
rect 262 133 279 137
rect 283 133 285 137
rect 262 132 285 133
rect 132 116 144 131
rect 148 131 169 132
rect 152 127 153 131
rect 157 128 169 131
rect 173 128 187 132
rect 191 128 205 132
rect 209 128 223 132
rect 227 128 241 132
rect 157 127 245 128
rect 148 126 245 127
rect 152 122 153 126
rect 157 122 245 126
rect 148 121 245 122
rect 262 128 279 132
rect 283 128 285 132
rect 262 127 285 128
rect 262 123 279 127
rect 283 123 285 127
rect 262 122 285 123
rect 262 118 279 122
rect 283 118 285 122
rect 262 117 285 118
rect 262 116 279 117
rect 0 112 2 116
rect 6 113 279 116
rect 283 113 285 117
rect 6 112 285 113
rect 0 108 137 112
rect 141 108 142 112
rect 146 108 147 112
rect 151 108 279 112
rect 283 108 285 112
rect 0 104 2 108
rect 6 107 285 108
rect 6 105 279 107
rect 6 104 142 105
rect 0 101 142 104
rect 146 101 150 105
rect 154 101 173 105
rect 177 101 185 105
rect 189 101 193 105
rect 197 101 211 105
rect 215 103 279 105
rect 283 103 285 107
rect 215 101 285 103
rect 0 100 285 101
rect 0 96 1 100
rect 5 99 285 100
rect 5 96 55 99
rect 0 95 55 96
rect 59 96 102 99
rect 59 95 80 96
rect 0 92 80 95
rect 84 95 102 96
rect 106 95 182 99
rect 186 97 213 99
rect 186 95 196 97
rect 84 93 196 95
rect 200 95 213 97
rect 217 95 232 99
rect 236 95 250 99
rect 254 95 274 99
rect 278 95 279 99
rect 283 95 285 99
rect 200 94 285 95
rect 200 93 213 94
rect 84 92 213 93
rect 0 91 196 92
rect 0 87 80 91
rect 84 90 196 91
rect 84 87 144 90
rect 0 86 144 87
rect 148 88 196 90
rect 200 90 213 92
rect 217 90 285 94
rect 200 88 285 90
rect 148 87 285 88
rect 148 86 196 87
rect 0 85 80 86
rect 0 81 1 85
rect 5 81 7 85
rect 11 81 23 85
rect 27 82 80 85
rect 84 85 196 86
rect 84 82 123 85
rect 27 81 123 82
rect 127 81 144 85
rect 148 83 196 85
rect 200 83 285 87
rect 148 82 285 83
rect 148 81 196 82
rect 0 78 196 81
rect 200 78 285 82
rect 0 77 285 78
rect 0 75 196 77
rect 0 71 8 75
rect 12 71 23 75
rect 27 71 46 75
rect 50 71 62 75
rect 66 74 139 75
rect 66 71 80 74
rect 0 70 80 71
rect 84 70 123 74
rect 127 71 139 74
rect 143 71 144 75
rect 148 71 167 75
rect 171 73 196 75
rect 200 73 285 77
rect 171 71 285 73
rect 127 70 285 71
rect 98 62 179 65
rect 0 57 1 61
rect 5 57 8 61
rect 12 58 13 61
rect 12 57 78 58
rect 82 57 285 58
rect 0 51 285 57
rect 0 47 7 51
rect 11 47 23 51
rect 27 50 285 51
rect 27 47 276 50
rect 0 46 276 47
rect 280 46 285 50
rect 0 44 132 46
rect 0 40 41 44
rect 45 42 132 44
rect 136 45 285 46
rect 136 44 276 45
rect 136 42 179 44
rect 45 41 179 42
rect 45 40 132 41
rect 0 37 132 40
rect 136 40 179 41
rect 183 41 276 44
rect 280 41 285 45
rect 183 40 285 41
rect 136 39 276 40
rect 136 37 179 39
rect 0 36 179 37
rect 0 32 132 36
rect 136 35 179 36
rect 183 36 276 39
rect 280 36 285 40
rect 183 35 285 36
rect 136 34 276 35
rect 136 32 179 34
rect 0 30 179 32
rect 183 31 276 34
rect 280 31 285 35
rect 183 30 285 31
rect 0 29 276 30
rect 0 25 179 29
rect 183 26 276 29
rect 280 26 285 30
rect 183 25 285 26
rect 0 24 276 25
rect 0 22 179 24
rect 0 18 1 22
rect 5 20 179 22
rect 183 23 276 24
rect 183 20 188 23
rect 5 19 188 20
rect 192 19 196 23
rect 200 19 204 23
rect 208 19 212 23
rect 216 19 220 23
rect 224 19 228 23
rect 232 19 236 23
rect 240 19 244 23
rect 248 19 252 23
rect 256 19 260 23
rect 264 21 276 23
rect 280 21 285 25
rect 264 20 285 21
rect 264 19 276 20
rect 5 18 276 19
rect 0 17 105 18
rect 0 13 1 17
rect 5 13 6 17
rect 10 13 23 17
rect 27 13 37 17
rect 41 13 47 17
rect 51 13 61 17
rect 65 13 81 17
rect 85 13 86 17
rect 90 14 105 17
rect 109 14 113 18
rect 117 14 121 18
rect 125 14 129 18
rect 133 14 137 18
rect 141 14 145 18
rect 149 14 153 18
rect 157 14 161 18
rect 165 14 174 18
rect 178 17 276 18
rect 178 14 192 17
rect 90 13 192 14
rect 196 13 200 17
rect 204 13 208 17
rect 212 13 216 17
rect 220 13 224 17
rect 228 13 232 17
rect 236 13 240 17
rect 244 13 248 17
rect 252 13 256 17
rect 260 13 264 17
rect 268 16 276 17
rect 280 16 285 20
rect 268 13 285 16
rect 0 10 285 13
rect 0 5 285 6
rect 0 1 7 5
rect 11 1 15 5
rect 19 1 23 5
rect 27 1 43 5
rect 47 1 80 5
rect 84 1 88 5
rect 92 1 105 5
rect 109 1 113 5
rect 117 1 121 5
rect 125 1 129 5
rect 133 1 137 5
rect 141 1 145 5
rect 149 1 153 5
rect 157 1 161 5
rect 165 1 179 5
rect 183 1 187 5
rect 191 1 195 5
rect 199 1 203 5
rect 207 1 211 5
rect 215 1 219 5
rect 223 1 227 5
rect 231 1 235 5
rect 239 1 243 5
rect 247 1 251 5
rect 255 1 259 5
rect 263 1 267 5
rect 271 1 275 5
rect 279 1 285 5
rect 0 0 285 1
<< ntransistor >>
rect 165 113 167 127
rect 175 111 177 127
rect 183 111 185 127
rect 193 111 195 127
rect 201 111 203 127
rect 211 111 213 127
rect 219 111 221 127
rect 229 111 231 127
rect 237 111 239 127
rect 247 111 249 127
rect 12 86 14 96
rect 20 86 22 96
rect 28 86 30 96
rect 36 86 38 96
rect 52 84 54 94
rect 60 84 62 94
rect 87 93 98 95
rect 112 84 114 96
rect 120 86 122 96
rect 128 86 130 96
rect 136 86 138 96
rect 156 84 158 96
rect 164 84 166 96
rect 172 84 174 96
<< ptransistor >>
rect 12 22 14 46
rect 20 22 22 46
rect 28 22 30 46
rect 36 22 38 46
rect 52 22 54 46
rect 60 22 62 46
rect 85 24 87 48
rect 106 24 108 46
rect 114 24 116 46
rect 122 24 124 46
rect 142 24 144 46
rect 150 24 152 46
rect 158 24 160 46
rect 166 24 168 48
rect 193 24 195 48
rect 201 24 203 48
rect 209 24 211 48
rect 217 24 219 48
rect 225 24 227 48
rect 233 24 235 48
rect 241 24 243 48
rect 249 24 251 48
rect 257 24 259 48
rect 265 24 267 48
<< polycontact >>
rect 162 108 166 112
rect 62 95 66 99
rect 38 81 42 85
rect 100 88 104 92
rect 104 81 108 85
rect 132 81 136 85
rect 182 81 186 85
rect 87 62 91 66
rect 104 62 108 66
rect 132 64 136 68
rect 165 64 169 68
rect 38 47 42 51
rect 62 47 66 51
rect 94 47 98 51
rect 108 47 112 51
rect 154 47 158 51
rect 179 47 183 51
rect 189 49 193 53
<< ndcontact >>
rect 1 142 5 314
rect 8 307 32 315
rect 11 294 27 302
rect 7 280 15 288
rect 20 277 28 293
rect 11 270 27 274
rect 6 259 14 263
rect 11 250 19 254
rect 7 241 15 245
rect 20 237 28 269
rect 11 227 27 235
rect 7 213 15 221
rect 20 209 28 225
rect 11 203 27 207
rect 7 193 15 197
rect 20 188 28 200
rect 11 179 27 187
rect 7 165 15 173
rect 10 156 18 160
rect 20 157 28 177
rect 10 151 18 155
rect 20 151 28 155
rect 34 203 42 315
rect 6 142 14 146
rect 34 143 42 171
rect 243 203 251 315
rect 254 307 278 315
rect 243 142 251 170
rect 258 294 274 302
rect 257 277 265 293
rect 270 280 278 288
rect 258 270 274 274
rect 257 236 265 268
rect 271 259 279 263
rect 266 250 274 254
rect 270 241 278 245
rect 258 227 274 235
rect 257 209 265 225
rect 270 213 278 221
rect 258 203 274 207
rect 257 188 265 200
rect 270 193 278 197
rect 258 179 274 187
rect 257 165 265 177
rect 270 165 278 173
rect 257 156 265 164
rect 267 156 275 160
rect 257 151 265 155
rect 267 151 275 155
rect 280 154 284 314
rect 252 142 256 146
rect 275 142 283 146
rect 12 109 28 129
rect 111 109 127 129
rect 160 116 164 127
rect 169 112 173 124
rect 178 112 182 124
rect 187 112 191 124
rect 196 112 200 124
rect 205 112 209 124
rect 214 112 218 124
rect 223 112 227 124
rect 232 112 236 124
rect 241 112 245 124
rect 250 112 254 124
rect 7 88 11 96
rect 15 88 19 96
rect 23 88 27 96
rect 31 88 35 96
rect 39 88 43 96
rect 47 87 51 94
rect 55 84 59 92
rect 63 84 67 92
rect 87 96 98 100
rect 87 88 95 92
rect 107 88 111 96
rect 115 84 119 96
rect 123 86 127 90
rect 131 88 135 96
rect 139 86 143 90
rect 151 84 155 96
rect 159 86 163 90
rect 167 92 171 96
rect 175 84 179 96
<< pdcontact >>
rect 214 64 222 80
rect 255 64 271 80
rect 7 22 11 46
rect 15 22 19 46
rect 23 22 27 46
rect 31 22 35 46
rect 39 22 43 40
rect 47 22 51 46
rect 55 22 59 46
rect 63 22 67 42
rect 80 24 84 48
rect 88 24 92 44
rect 101 25 105 45
rect 109 24 113 36
rect 117 32 121 44
rect 125 25 129 45
rect 137 30 141 46
rect 145 24 149 36
rect 153 32 157 44
rect 161 25 165 45
rect 174 25 178 41
rect 188 24 192 44
rect 196 28 200 48
rect 204 24 208 48
rect 212 28 216 48
rect 220 24 224 48
rect 228 28 232 48
rect 236 24 240 48
rect 244 28 248 48
rect 252 24 256 48
rect 260 28 264 48
rect 268 24 272 48
<< m2contact >>
rect 2 132 6 136
rect 2 124 6 128
rect 2 112 6 116
rect 2 104 6 108
rect 11 135 15 139
rect 133 131 137 135
rect 138 131 142 135
rect 148 127 152 131
rect 153 127 157 131
rect 148 122 152 126
rect 153 122 157 126
rect 169 128 173 132
rect 1 96 5 100
rect 1 81 5 85
rect 7 81 11 85
rect 8 71 12 75
rect 8 66 12 70
rect 55 95 59 99
rect 137 108 141 112
rect 142 108 146 112
rect 147 108 151 112
rect 142 101 146 105
rect 150 101 154 105
rect 23 81 27 85
rect 23 71 27 75
rect 23 66 27 70
rect 1 57 5 61
rect 8 57 12 61
rect 7 47 11 51
rect 23 47 27 51
rect 46 71 50 75
rect 46 66 50 70
rect 62 71 66 75
rect 62 66 66 70
rect 1 18 5 22
rect 1 13 5 17
rect 6 13 10 17
rect 23 13 27 17
rect 80 92 84 96
rect 102 95 106 99
rect 187 128 191 132
rect 205 128 209 132
rect 173 101 177 105
rect 185 101 189 105
rect 193 101 197 105
rect 80 87 84 91
rect 80 82 84 86
rect 80 70 84 74
rect 78 57 82 61
rect 41 40 45 44
rect 7 1 11 5
rect 15 1 19 5
rect 23 1 27 5
rect 37 13 41 17
rect 47 13 51 17
rect 43 1 47 5
rect 61 13 65 17
rect 94 62 98 66
rect 144 86 148 90
rect 81 13 85 17
rect 86 13 90 17
rect 80 1 84 5
rect 88 1 92 5
rect 123 81 127 85
rect 123 70 127 74
rect 144 81 148 85
rect 182 95 186 99
rect 196 93 200 97
rect 139 71 143 75
rect 144 71 148 75
rect 167 71 171 75
rect 179 62 183 66
rect 132 42 136 46
rect 132 37 136 41
rect 132 32 136 36
rect 105 14 109 18
rect 113 14 117 18
rect 121 14 125 18
rect 129 14 133 18
rect 137 14 141 18
rect 145 14 149 18
rect 153 14 157 18
rect 161 14 165 18
rect 105 1 109 5
rect 113 1 117 5
rect 121 1 125 5
rect 129 1 133 5
rect 137 1 141 5
rect 145 1 149 5
rect 153 1 157 5
rect 161 1 165 5
rect 196 88 200 92
rect 196 83 200 87
rect 196 78 200 82
rect 223 128 227 132
rect 211 101 215 105
rect 213 95 217 99
rect 213 90 217 94
rect 232 95 236 99
rect 241 128 245 132
rect 250 95 254 99
rect 279 133 283 137
rect 279 128 283 132
rect 279 123 283 127
rect 279 118 283 122
rect 279 113 283 117
rect 279 108 283 112
rect 279 103 283 107
rect 274 95 278 99
rect 279 95 283 99
rect 196 73 200 77
rect 179 40 183 44
rect 179 35 183 39
rect 179 30 183 34
rect 179 25 183 29
rect 179 20 183 24
rect 188 19 192 23
rect 196 19 200 23
rect 204 19 208 23
rect 212 19 216 23
rect 220 19 224 23
rect 228 19 232 23
rect 236 19 240 23
rect 244 19 248 23
rect 252 19 256 23
rect 260 19 264 23
rect 276 46 280 50
rect 276 41 280 45
rect 276 36 280 40
rect 276 31 280 35
rect 276 26 280 30
rect 276 21 280 25
rect 174 14 178 18
rect 192 13 196 17
rect 200 13 204 17
rect 208 13 212 17
rect 216 13 220 17
rect 224 13 228 17
rect 232 13 236 17
rect 240 13 244 17
rect 248 13 252 17
rect 256 13 260 17
rect 264 13 268 17
rect 276 16 280 20
rect 179 1 183 5
rect 187 1 191 5
rect 195 1 199 5
rect 203 1 207 5
rect 211 1 215 5
rect 219 1 223 5
rect 227 1 231 5
rect 235 1 239 5
rect 243 1 247 5
rect 251 1 255 5
rect 259 1 263 5
rect 267 1 271 5
rect 275 1 279 5
<< psubstratepcontact >>
rect 2 136 6 140
rect 7 135 11 139
rect 33 135 141 139
rect 159 135 163 139
rect 178 135 182 139
rect 196 135 200 139
rect 214 135 218 139
rect 232 135 236 139
rect 250 135 254 139
rect 2 128 6 132
rect 2 116 6 124
rect 2 108 6 112
rect 3 100 27 104
rect 29 100 33 104
rect 34 100 42 104
rect 3 87 7 95
rect 43 88 47 104
rect 49 100 53 104
rect 55 100 59 104
rect 78 100 126 104
rect 138 101 142 105
rect 146 101 150 105
rect 154 101 158 105
rect 169 101 173 105
rect 177 101 185 105
rect 189 101 193 105
rect 197 101 201 105
rect 215 101 219 105
rect 232 102 236 106
rect 250 102 254 106
rect 275 100 279 140
rect 189 95 193 99
rect 23 76 27 80
rect 46 76 50 80
rect 62 76 66 80
rect 80 76 84 80
rect 123 76 127 80
rect 139 76 143 80
rect 144 76 148 80
rect 150 76 154 80
rect 167 76 171 80
rect 3 1 7 5
rect 11 1 15 5
rect 19 1 23 5
rect 39 1 43 5
rect 47 1 51 5
rect 76 1 80 5
rect 84 1 88 5
rect 101 1 105 5
rect 109 1 113 5
rect 117 1 121 5
rect 125 1 129 5
rect 133 1 137 5
rect 141 1 145 5
rect 149 1 153 5
rect 157 1 161 5
rect 175 1 179 5
rect 183 1 187 5
rect 191 1 195 5
rect 199 1 203 5
rect 207 1 211 5
rect 215 1 219 5
rect 223 1 227 5
rect 231 1 235 5
rect 239 1 243 5
rect 247 1 251 5
rect 255 1 259 5
rect 263 1 267 5
rect 271 1 275 5
<< nsubstratencontact >>
rect 1 52 5 56
rect 7 52 11 56
rect 23 52 27 56
rect 47 52 51 56
rect 78 52 82 56
rect 3 22 7 46
rect 43 20 47 40
rect 11 13 23 17
rect 42 12 46 16
rect 76 12 80 48
rect 133 50 137 54
rect 147 52 151 56
rect 204 54 208 58
rect 220 54 224 58
rect 236 54 240 58
rect 268 54 272 58
rect 276 52 284 88
rect 184 24 188 44
rect 272 21 276 49
rect 280 18 284 50
rect 101 14 105 18
rect 109 14 113 18
rect 117 14 121 18
rect 125 14 129 18
rect 133 14 137 18
rect 141 14 145 18
rect 149 14 153 18
rect 157 14 161 18
rect 184 14 192 18
rect 196 14 200 18
rect 204 14 208 18
rect 212 14 216 18
rect 220 14 224 18
rect 228 14 232 18
rect 236 14 240 18
rect 244 14 248 18
rect 252 14 256 18
rect 260 14 264 18
rect 268 14 276 18
<< psubstratepdiff >>
rect 0 140 285 141
rect 0 136 2 140
rect 6 139 275 140
rect 6 136 7 139
rect 0 135 7 136
rect 11 135 33 139
rect 141 135 159 139
rect 163 135 178 139
rect 182 135 196 139
rect 200 135 214 139
rect 218 135 232 139
rect 236 135 250 139
rect 254 135 275 139
rect 0 133 275 135
rect 0 132 8 133
rect 0 128 2 132
rect 6 128 8 132
rect 0 124 8 128
rect 0 116 2 124
rect 6 116 8 124
rect 0 112 8 116
rect 0 108 2 112
rect 6 108 8 112
rect 0 105 8 108
rect 131 107 160 133
rect 254 107 275 133
rect 131 106 275 107
rect 131 105 232 106
rect 0 104 138 105
rect 0 100 3 104
rect 27 100 29 104
rect 33 100 34 104
rect 42 100 43 104
rect 0 96 6 100
rect 0 95 7 96
rect 0 87 3 95
rect 0 86 7 87
rect 47 100 49 104
rect 53 100 55 104
rect 59 100 78 104
rect 126 101 138 104
rect 142 101 146 105
rect 150 101 154 105
rect 158 101 169 105
rect 173 101 177 105
rect 185 101 189 105
rect 193 101 197 105
rect 201 101 215 105
rect 219 102 232 105
rect 236 102 250 106
rect 254 102 275 106
rect 219 101 275 102
rect 126 100 275 101
rect 279 100 285 140
rect 0 80 6 86
rect 43 80 47 88
rect 67 80 74 100
rect 187 99 195 100
rect 187 95 189 99
rect 193 95 195 99
rect 187 80 195 95
rect 0 76 23 80
rect 27 76 46 80
rect 50 76 62 80
rect 66 76 80 80
rect 84 76 123 80
rect 127 76 139 80
rect 143 76 144 80
rect 148 76 150 80
rect 154 76 167 80
rect 171 76 195 80
rect 0 5 285 6
rect 0 1 3 5
rect 7 1 11 5
rect 15 1 19 5
rect 23 1 39 5
rect 43 1 47 5
rect 51 1 76 5
rect 80 1 84 5
rect 88 1 101 5
rect 105 1 109 5
rect 113 1 117 5
rect 121 1 125 5
rect 129 1 133 5
rect 137 1 141 5
rect 145 1 149 5
rect 153 1 157 5
rect 161 1 175 5
rect 179 1 183 5
rect 187 1 191 5
rect 195 1 199 5
rect 203 1 207 5
rect 211 1 215 5
rect 219 1 223 5
rect 227 1 231 5
rect 235 1 239 5
rect 243 1 247 5
rect 251 1 255 5
rect 259 1 263 5
rect 267 1 271 5
rect 275 1 285 5
rect 0 0 285 1
<< nsubstratendiff >>
rect 204 88 285 89
rect 204 85 276 88
rect 204 59 210 85
rect 275 59 276 85
rect 184 58 276 59
rect 184 56 204 58
rect 0 52 1 56
rect 5 52 7 56
rect 11 52 23 56
rect 27 52 47 56
rect 51 52 78 56
rect 82 54 147 56
rect 82 52 133 54
rect 0 46 6 52
rect 0 22 3 46
rect 43 40 47 52
rect 67 48 80 52
rect 0 18 7 22
rect 43 18 47 20
rect 67 18 76 48
rect 0 17 76 18
rect 0 13 11 17
rect 23 16 76 17
rect 23 13 42 16
rect 0 12 42 13
rect 46 12 76 16
rect 131 50 133 52
rect 137 52 147 54
rect 151 54 204 56
rect 208 54 220 58
rect 224 54 236 58
rect 240 54 268 58
rect 151 52 188 54
rect 137 50 141 52
rect 184 46 188 52
rect 272 52 276 58
rect 284 52 285 88
rect 272 50 285 52
rect 272 49 280 50
rect 178 44 188 46
rect 178 24 184 44
rect 174 20 187 24
rect 80 18 187 20
rect 276 21 280 49
rect 272 18 280 21
rect 284 18 285 50
rect 80 14 101 18
rect 105 14 109 18
rect 113 14 117 18
rect 121 14 125 18
rect 129 14 133 18
rect 137 14 141 18
rect 145 14 149 18
rect 153 14 157 18
rect 161 14 184 18
rect 192 14 196 18
rect 200 14 204 18
rect 208 14 212 18
rect 216 14 220 18
rect 224 14 228 18
rect 232 14 236 18
rect 240 14 244 18
rect 248 14 252 18
rect 256 14 260 18
rect 264 14 268 18
rect 276 14 285 18
rect 80 12 285 14
<< pad >>
rect 72 173 214 315
<< glass >>
rect 78 179 208 309
<< labels >>
rlabel metal1 96 0 96 0 8 EN
rlabel metal1 169 0 169 0 8 OUT
rlabel metal2 93 22 93 22 6 Vdd
rlabel pdcontact 147 30 147 30 6 P
rlabel polysilicon 167 49 167 49 6 EN
rlabel polysilicon 149 48 149 48 6 OUT
rlabel polysilicon 123 48 123 48 6 ENB
rlabel pdcontact 103 28 103 28 6 N
rlabel metal2 92 84 92 84 6 GND
rlabel ndcontact 116 90 116 90 6 N
rlabel ndcontact 133 90 133 90 6 N
rlabel polysilicon 121 85 121 85 6 OUT
rlabel polysilicon 113 83 113 83 6 ENB
rlabel ndcontact 161 88 161 88 6 P
rlabel polysilicon 165 82 165 82 6 EN
rlabel space 0 320 0 320 4 sllu_1988
rlabel metal1 32 0 32 0 8 IN
rlabel space 285 320 285 320 6 mosis_tinychip
rlabel metal1 143 234 143 234 6 pad
rlabel metal1 71 0 71 0 8 in_unbuf
rlabel space 147 153 147 153 6 1989
rlabel space 147 155 147 155 6 MOSIS
rlabel space 147 157 147 157 6 Shih-Lien_Lu
rlabel metal2 0 70 0 70 4 {w}tiny12_t
rlabel nsubstratendiff 285 70 285 70 6 {e}tiny12_t
rlabel nsubstratendiff 285 58 285 58 6 {e}tiny12_b
rlabel metal2 0 58 0 58 4 {w}tiny12_b
rlabel metal1 56 0 56 0 8 INb
rlabel psubstratepdiff 0 100 0 100 4 {w}tiny12_L
rlabel psubstratepdiff 285 100 285 100 6 {e}tiny12_R
<< end >>
