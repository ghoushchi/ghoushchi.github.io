magic
tech scmos
timestamp 951255912
<< metal2 >>
rect 12 180 16 210
rect 12 116 16 146
rect 12 54 16 84
use memtile memtile_3
timestamp 951255912
transform 1 0 95 0 1 192
box -95 -1 451 69
use memtile memtile_2
timestamp 951255912
transform 1 0 95 0 1 128
box -95 -1 451 69
use memtile memtile_1
timestamp 951255912
transform 1 0 95 0 1 64
box -95 -1 451 69
use memtile memtile_0
timestamp 951255912
transform 1 0 95 0 1 0
box -95 -1 451 69
<< end >>
