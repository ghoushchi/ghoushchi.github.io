magic
tech scmos
timestamp 951209823
<< nwell >>
rect 77 39 115 71
<< polysilicon >>
rect 89 64 108 66
rect 89 63 91 64
rect 89 53 91 55
rect 97 51 99 53
rect 89 49 91 51
rect 89 39 91 41
rect 85 37 91 39
rect 85 23 87 37
rect 97 30 99 41
rect 98 26 99 30
rect 89 23 91 25
rect 97 23 99 26
rect 97 16 99 18
rect 85 13 87 15
rect 89 14 91 15
rect 89 12 108 14
<< ndiffusion >>
rect 84 15 85 23
rect 87 15 89 23
rect 91 15 92 23
rect 96 18 97 23
rect 99 18 100 23
<< pdiffusion >>
rect 88 55 89 63
rect 91 55 92 63
rect 88 41 89 49
rect 91 41 92 49
rect 96 41 97 51
rect 99 41 100 51
<< metal1 >>
rect 89 67 92 71
rect 92 63 96 67
rect 84 49 88 55
rect 80 29 84 49
rect 92 51 96 55
rect 108 66 112 71
rect 91 33 92 37
rect 80 26 94 29
rect 101 28 104 41
rect 80 23 84 26
rect 101 23 104 24
rect 92 11 96 15
rect 89 7 92 11
rect 108 16 112 62
rect 108 7 112 12
<< metal2 >>
rect 77 67 92 71
rect 96 67 112 71
rect 77 66 112 67
rect 80 33 92 37
rect 77 29 84 33
rect 105 24 108 28
rect 77 11 112 12
rect 77 7 92 11
rect 96 7 112 11
<< ntransistor >>
rect 85 15 87 23
rect 89 15 91 23
rect 97 18 99 23
<< ptransistor >>
rect 89 55 91 63
rect 89 41 91 49
rect 97 41 99 51
<< polycontact >>
rect 108 62 112 66
rect 87 33 91 37
rect 94 26 98 30
rect 108 12 112 16
<< ndcontact >>
rect 80 15 84 23
rect 92 15 96 23
rect 100 18 104 23
<< pdcontact >>
rect 84 55 88 63
rect 92 55 96 63
rect 84 41 88 49
rect 92 41 96 51
rect 100 41 104 51
<< m2contact >>
rect 92 67 96 71
rect 92 33 96 37
rect 101 24 105 28
rect 92 7 96 11
<< psubstratepcontact >>
rect 82 7 89 11
<< nsubstratencontact >>
rect 82 67 89 71
<< labels >>
rlabel metal2 100 9 100 9 5 Gnd
rlabel metal2 101 69 101 69 1 Vdd
rlabel metal2 80 31 80 31 7 FromMux
rlabel metal2 106 26 106 26 3 ToAdd
rlabel metal1 110 9 110 9 5 PixBit
<< end >>
