magic
tech scmos
timestamp 951308881
<< nwell >>
rect -10 -10 14 22
<< polysilicon >>
rect -2 46 0 48
rect 6 46 8 48
rect -2 34 0 36
rect 6 34 8 36
rect -2 32 8 34
rect -3 28 0 32
rect -2 18 0 28
rect 6 18 8 32
rect -2 -4 0 -2
rect 6 -4 8 -2
<< ndiffusion >>
rect -3 36 -2 46
rect 0 36 1 46
rect 5 36 6 46
rect 8 36 9 46
<< pdiffusion >>
rect -3 -2 -2 18
rect 0 -2 1 18
rect 5 -2 6 18
rect 8 -2 9 18
<< metal1 >>
rect -7 50 -1 54
rect 7 50 13 54
rect -7 46 -3 50
rect 9 46 13 50
rect -7 27 -3 28
rect 1 27 5 36
rect 1 23 9 27
rect 1 18 5 23
rect -7 -6 -3 -2
rect 9 -6 13 -2
rect -7 -10 -1 -6
rect 7 -10 13 -6
<< ntransistor >>
rect -2 36 0 46
rect 6 36 8 46
<< ptransistor >>
rect -2 -2 0 18
rect 6 -2 8 18
<< polycontact >>
rect -7 28 -3 32
<< ndcontact >>
rect -7 36 -3 46
rect 1 36 5 46
rect 9 36 13 46
<< pdcontact >>
rect -7 -2 -3 18
rect 1 -2 5 18
rect 9 -2 13 18
<< m2contact >>
rect -7 23 -3 27
rect 9 23 13 27
<< psubstratepcontact >>
rect -1 50 7 54
<< nsubstratencontact >>
rect -1 -10 7 -6
<< labels >>
rlabel m2contact -5 25 -5 25 3 In
rlabel psubstratepcontact 3 52 3 52 5 Gnd
rlabel nsubstratencontact 3 -8 3 -8 1 Vdd
rlabel m2contact 11 25 11 25 7 Out
<< end >>
