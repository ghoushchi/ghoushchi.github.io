magic
tech scmos
timestamp 951112323
<< metal1 >>
rect 11 79 14 87
rect 18 79 21 83
rect 119 79 122 87
rect 126 79 129 83
rect 167 20 172 127
rect 63 -99 70 -96
rect 167 -100 172 14
rect 175 -40 180 74
rect 175 -105 180 -46
<< metal2 >>
rect 12 127 167 132
rect 11 95 15 99
rect 119 95 124 99
rect 27 74 32 79
rect 167 74 175 79
rect 3 40 9 44
rect 4 -10 10 -6
rect 167 -46 175 -40
rect 4 -80 9 -76
rect 28 -105 35 -100
<< m2contact >>
rect 167 127 172 132
rect 11 87 15 91
rect 119 87 123 91
rect 167 14 172 20
rect 167 -105 172 -100
rect 175 74 180 79
rect 175 -46 180 -40
use inverters inverters_1
timestamp 951078626
transform 1 0 49 0 1 87
box -37 -12 2 45
use inverters inverters_0
timestamp 951078626
transform 1 0 157 0 1 87
box -37 -12 2 45
use SetCell SetCell_0
timestamp 951088720
transform 1 0 20 0 1 18
box -17 -3 147 61
use ResetCell ResetCell_0
timestamp 951088720
transform 1 0 25 0 -1 6
box -21 -13 142 51
use ResetCellflip ResetCellflip_0
timestamp 951112323
transform 1 0 -5 0 1 -192
box 9 87 172 151
<< labels >>
rlabel metal2 30 76 30 76 5 Vdd
rlabel metal2 32 -103 32 -103 1 Gnd
rlabel metal2 4 42 4 42 3 kernelCounterOut2_s1
rlabel metal2 5 -9 5 -9 3 kernelCounterOut1_s1
rlabel metal2 5 -79 5 -79 3 kernelCounterOut0_s1
rlabel metal2 12 97 12 97 1 c3_Phi2_q2
rlabel metal2 120 97 120 97 1 Phi1
<< end >>
