magic
tech scmos
timestamp 950486748
<< polysilicon >>
rect 244 114 259 150
rect 205 100 297 114
rect 244 62 259 100
<< metal1 >>
rect 162 167 330 335
rect 3 130 126 131
rect 3 126 4 130
rect 8 126 9 130
rect 13 126 14 130
rect 18 126 126 130
rect 3 125 126 126
rect 3 121 4 125
rect 8 121 9 125
rect 13 121 14 125
rect 18 121 126 125
rect 3 120 126 121
rect 3 116 4 120
rect 8 116 9 120
rect 13 116 14 120
rect 18 116 126 120
rect 3 115 126 116
rect 3 111 4 115
rect 8 111 9 115
rect 13 111 14 115
rect 18 111 126 115
rect 3 110 126 111
rect 3 106 4 110
rect 8 106 9 110
rect 13 106 14 110
rect 18 106 126 110
rect 3 105 126 106
rect 3 101 4 105
rect 8 101 9 105
rect 13 101 14 105
rect 18 101 126 105
rect 3 100 126 101
rect 3 96 4 100
rect 8 96 9 100
rect 13 96 14 100
rect 18 96 126 100
rect 3 95 126 96
rect 3 91 4 95
rect 8 91 9 95
rect 13 91 14 95
rect 18 91 126 95
rect 3 90 126 91
rect 3 86 4 90
rect 8 86 9 90
rect 13 86 14 90
rect 18 86 126 90
rect 3 85 126 86
rect 7 83 126 85
rect 10 21 15 83
rect 20 55 55 60
rect 20 47 21 55
rect 29 54 55 55
rect 29 47 33 54
rect 20 38 33 47
rect 7 20 16 21
rect 15 16 16 20
rect 11 15 16 16
rect 15 7 16 15
rect 29 10 33 38
rect 41 46 55 54
rect 41 42 45 46
rect 49 42 50 46
rect 54 42 55 46
rect 41 41 55 42
rect 41 37 45 41
rect 49 37 50 41
rect 54 37 55 41
rect 41 10 55 37
rect 29 7 55 10
rect 75 13 126 83
rect 75 9 81 13
rect 85 9 86 13
rect 90 9 91 13
rect 95 9 96 13
rect 100 9 101 13
rect 105 9 106 13
rect 110 9 111 13
rect 115 9 116 13
rect 120 9 121 13
rect 125 9 126 13
rect 75 8 126 9
rect 75 6 81 8
rect 80 4 81 6
rect 85 4 86 8
rect 90 4 91 8
rect 95 4 96 8
rect 100 4 101 8
rect 105 4 106 8
rect 110 4 111 8
rect 115 4 116 8
rect 120 4 121 8
rect 125 4 126 8
<< metal2 >>
rect 27 330 329 334
rect 27 172 167 330
rect 325 172 329 330
rect 27 168 329 172
rect 0 130 18 131
rect 0 126 4 130
rect 8 126 9 130
rect 13 126 14 130
rect 0 125 18 126
rect 0 121 4 125
rect 8 121 9 125
rect 13 121 14 125
rect 0 120 18 121
rect 0 116 4 120
rect 8 116 9 120
rect 13 116 14 120
rect 0 115 18 116
rect 0 111 4 115
rect 8 111 9 115
rect 13 111 14 115
rect 0 110 18 111
rect 0 106 4 110
rect 8 106 9 110
rect 13 106 14 110
rect 0 105 18 106
rect 0 101 4 105
rect 8 101 9 105
rect 13 101 14 105
rect 0 100 18 101
rect 0 96 4 100
rect 8 96 9 100
rect 13 96 14 100
rect 0 95 18 96
rect 0 91 4 95
rect 8 91 9 95
rect 13 91 14 95
rect 0 90 18 91
rect 0 86 4 90
rect 8 86 9 90
rect 13 86 14 90
rect 0 85 18 86
rect 27 73 163 168
rect 0 46 163 73
rect 0 42 45 46
rect 49 42 50 46
rect 54 42 163 46
rect 0 41 163 42
rect 0 37 45 41
rect 49 37 50 41
rect 54 37 163 41
rect 0 25 163 37
rect 20 22 163 25
rect 0 20 16 21
rect 0 16 3 20
rect 7 16 11 20
rect 15 16 16 20
rect 0 15 16 16
rect 10 11 16 15
rect 10 7 11 11
rect 15 7 16 11
rect 10 0 16 7
rect 20 0 68 22
rect 80 9 81 13
rect 85 9 86 13
rect 90 9 91 13
rect 95 9 96 13
rect 100 9 101 13
rect 105 9 106 13
rect 110 9 111 13
rect 115 9 116 13
rect 120 9 121 13
rect 125 9 126 13
rect 80 8 126 9
rect 80 4 81 8
rect 85 4 86 8
rect 90 4 91 8
rect 95 4 96 8
rect 100 4 101 8
rect 105 4 106 8
rect 110 4 111 8
rect 115 4 116 8
rect 120 4 121 8
rect 125 4 126 8
rect 80 0 126 4
<< m2contact >>
rect 4 126 8 130
rect 9 126 13 130
rect 14 126 18 130
rect 4 121 8 125
rect 9 121 13 125
rect 14 121 18 125
rect 4 116 8 120
rect 9 116 13 120
rect 14 116 18 120
rect 4 111 8 115
rect 9 111 13 115
rect 14 111 18 115
rect 4 106 8 110
rect 9 106 13 110
rect 14 106 18 110
rect 4 101 8 105
rect 9 101 13 105
rect 14 101 18 105
rect 4 96 8 100
rect 9 96 13 100
rect 14 96 18 100
rect 4 91 8 95
rect 9 91 13 95
rect 14 91 18 95
rect 4 86 8 90
rect 9 86 13 90
rect 14 86 18 90
rect 3 16 7 20
rect 11 16 15 20
rect 11 7 15 11
rect 45 42 49 46
rect 50 42 54 46
rect 45 37 49 41
rect 50 37 54 41
rect 81 9 85 13
rect 86 9 90 13
rect 91 9 95 13
rect 96 9 100 13
rect 101 9 105 13
rect 106 9 110 13
rect 111 9 115 13
rect 116 9 120 13
rect 121 9 125 13
rect 81 4 85 8
rect 86 4 90 8
rect 91 4 95 8
rect 96 4 100 8
rect 101 4 105 8
rect 106 4 110 8
rect 111 4 115 8
rect 116 4 120 8
rect 121 4 125 8
<< psubstratepcontact >>
rect 7 16 11 20
rect 11 11 15 15
<< nsubstratencontact >>
rect 21 47 29 55
rect 33 10 41 54
<< psubstratepdiff >>
rect 0 20 16 21
rect 0 16 7 20
rect 11 16 16 20
rect 0 15 16 16
rect 10 11 11 15
rect 15 11 16 15
rect 10 0 16 11
<< nsubstratendiff >>
rect 0 55 66 71
rect 0 47 21 55
rect 29 54 66 55
rect 29 47 33 54
rect 0 27 33 47
rect 22 10 33 27
rect 41 10 66 54
rect 22 0 66 10
<< pad >>
rect 167 172 325 330
<< glass >>
rect 173 178 319 324
<< labels >>
rlabel metal2 44 57 44 57 6 Vdd
rlabel metal1 330 335 330 335 6 sllu
rlabel space 330 0 330 0 8 sllu_1988
rlabel space 0 335 0 335 4 sllu_1988
rlabel metal2 0 73 0 73 4 {w}tiny12_b
rlabel metal2 0 85 0 85 4 {w}tiny12_t
rlabel metal2 68 0 68 0 8 {s}tiny12_b
rlabel metal2 80 0 80 0 8 {s}tiny12_t
rlabel metal2 110 0 110 0 8 {s}*
rlabel metal2 0 115 0 115 4 {w}*
<< end >>
