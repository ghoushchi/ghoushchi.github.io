magic
tech scmos
timestamp 951288779
<< nwell >>
rect 9 -7 30 29
<< polysilicon >>
rect -6 22 -3 24
rect 2 22 12 24
rect 22 22 24 24
rect -6 5 -4 22
rect 4 13 8 15
rect 4 11 20 13
rect 18 5 20 11
rect -6 3 -3 5
rect 2 3 4 5
rect 10 3 12 5
rect 17 3 20 5
<< ndiffusion >>
rect -3 24 2 25
rect -3 21 2 22
rect -3 5 2 6
rect -3 2 2 3
<< pdiffusion >>
rect 12 24 22 25
rect 12 21 22 22
rect 12 5 17 6
rect 12 2 17 3
<< metal1 >>
rect -67 -7 -63 29
rect -60 -7 -56 29
rect -53 -7 -49 29
rect -46 -7 -42 29
rect -39 -7 -35 29
rect -32 -7 -28 29
rect -25 -7 -21 29
rect -18 -7 -14 29
rect -7 25 -3 29
rect 22 25 30 29
rect -11 -7 -6 25
rect 2 19 12 21
rect 2 17 4 19
rect 8 18 12 19
rect 25 11 30 25
rect 2 6 5 9
rect 9 6 12 9
rect 2 -2 5 1
rect 9 -2 12 1
rect 25 -7 30 7
<< metal2 >>
rect -70 9 9 13
rect 9 -3 34 1
<< ntransistor >>
rect -3 22 2 24
rect -3 3 2 5
<< ptransistor >>
rect 12 22 22 24
rect 12 3 17 5
<< polycontact >>
rect 4 15 8 19
<< ndcontact >>
rect -3 25 2 29
rect -3 17 2 21
rect -3 6 2 10
rect -3 -2 2 2
<< pdcontact >>
rect 12 25 22 29
rect 12 17 22 21
rect 12 6 17 10
rect 12 -2 17 2
<< m2contact >>
rect 5 5 9 9
rect 5 -3 9 1
rect 34 -3 38 1
<< psubstratepcontact >>
rect -11 25 -7 29
<< nsubstratencontact >>
rect 25 7 30 11
<< labels >>
rlabel psubstratepcontact -9 21 -9 21 1 Gnd
rlabel m2contact 7 -1 7 -1 1 out
rlabel m2contact 7 7 7 7 1 in
rlabel metal1 27 20 27 20 7 Vdd
<< end >>
