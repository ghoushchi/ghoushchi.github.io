magic
tech scmos
timestamp 943334529
<< pwell >>
rect -22 -2 63 34
<< nwell >>
rect -22 34 63 62
<< polysilicon >>
rect -7 57 -5 59
rect 9 57 11 59
rect 46 57 48 59
rect 50 57 52 59
rect 54 57 56 59
rect -7 48 -5 49
rect -12 46 -5 48
rect 9 48 11 49
rect 9 46 33 48
rect -12 34 -10 46
rect 46 42 48 45
rect 0 40 48 42
rect -12 32 -5 34
rect -7 7 -5 32
rect 9 7 11 40
rect 50 36 52 45
rect 46 34 52 36
rect 46 33 48 34
rect 45 29 48 33
rect 37 20 40 24
rect 38 17 40 20
rect 46 17 48 29
rect 54 25 56 45
rect 54 21 57 25
rect 54 17 56 21
rect 38 11 40 13
rect 46 11 48 13
rect 54 11 56 13
rect -7 1 -5 3
rect 9 1 11 3
<< ndiffusion >>
rect 37 13 38 17
rect 40 13 41 17
rect 45 13 46 17
rect 48 13 49 17
rect 53 13 54 17
rect 56 13 57 17
rect -8 3 -7 7
rect -5 3 -4 7
rect 8 3 9 7
rect 11 3 12 7
<< pdiffusion >>
rect -8 49 -7 57
rect -5 49 -4 57
rect 8 49 9 57
rect 11 49 12 57
rect 45 45 46 57
rect 48 45 50 57
rect 52 45 54 57
rect 56 45 57 57
<< metal1 >>
rect -19 54 -15 62
rect -19 24 -15 50
rect -12 57 -8 58
rect -4 42 0 49
rect -19 20 -11 24
rect -19 -2 -15 20
rect -12 7 -8 11
rect -4 7 0 38
rect 4 30 8 49
rect 4 7 8 26
rect 12 22 16 49
rect 12 7 16 18
rect 19 30 23 62
rect -12 2 -8 3
rect 19 -2 23 26
rect 26 38 30 62
rect 37 58 41 62
rect 41 57 45 58
rect 26 -2 30 34
rect 33 49 37 50
rect 33 24 37 45
rect 57 38 61 45
rect 41 33 45 34
rect 49 34 57 38
rect 49 22 53 34
rect 57 25 61 26
rect 49 17 53 18
rect 33 2 37 13
rect 41 10 45 13
rect 57 10 61 13
rect 41 6 61 10
<< metal2 >>
rect -22 58 -12 62
rect -8 58 41 62
rect 45 58 63 62
rect -15 50 33 54
rect -22 42 63 46
rect 30 34 41 38
rect 61 34 63 38
rect -22 26 4 30
rect 23 26 57 30
rect 16 18 49 22
rect -22 10 62 14
rect -22 -2 -12 2
rect -8 -2 33 2
rect 37 -2 63 2
<< ntransistor >>
rect 38 13 40 17
rect 46 13 48 17
rect 54 13 56 17
rect -7 3 -5 7
rect 9 3 11 7
<< ptransistor >>
rect -7 49 -5 57
rect 9 49 11 57
rect 46 45 48 57
rect 50 45 52 57
rect 54 45 56 57
<< polycontact >>
rect 33 45 37 49
rect -4 38 0 42
rect -11 20 -7 24
rect 41 29 45 33
rect 33 20 37 24
rect 57 21 61 25
<< ndcontact >>
rect 33 13 37 17
rect 41 13 45 17
rect 49 13 53 17
rect 57 13 61 17
rect -12 3 -8 7
rect -4 3 0 7
rect 4 3 8 7
rect 12 3 16 7
<< pdcontact >>
rect -12 49 -8 57
rect -4 49 0 57
rect 4 49 8 57
rect 12 49 16 57
rect 41 45 45 57
rect 57 45 61 57
<< m2contact >>
rect -19 50 -15 54
rect -12 58 -8 62
rect 4 26 8 30
rect 12 18 16 22
rect 19 26 23 30
rect -12 -2 -8 2
rect 41 58 45 62
rect 26 34 30 38
rect 33 50 37 54
rect 41 34 45 38
rect 57 34 61 38
rect 49 18 53 22
rect 57 26 61 30
rect 33 -2 37 2
<< psubstratepcontact >>
rect -12 11 -8 15
<< nsubstratencontact >>
rect 33 58 37 62
<< labels >>
rlabel metal2 60 0 60 0 3 Gnd
rlabel metal2 60 60 60 60 3 Vdd
rlabel metal2 -20 28 -20 28 7 in
rlabel metal1 -17 0 -17 0 7 reset_sr_s2
rlabel metal1 21 -1 21 -1 6 bits_s2[0]
rlabel metal1 28 -1 28 -1 4 coeff_en_b_s2
rlabel metal2 62 36 62 36 3 out
<< end >>
