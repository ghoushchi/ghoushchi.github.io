magic
tech scmos
timestamp 951985653
<< metal1 >>
rect 610 686 630 690
rect 610 679 622 683
rect 606 643 614 647
rect 34 524 74 528
rect 3 482 46 483
rect 0 479 46 482
rect 0 478 6 479
rect 3 386 46 389
rect 0 385 46 386
rect 0 382 6 385
rect 34 340 73 344
rect 89 262 101 266
rect 105 262 640 266
rect 155 254 640 258
rect 225 246 640 250
rect 275 238 640 242
rect 345 230 640 234
rect 395 222 640 226
rect 465 214 640 218
rect 515 206 640 210
rect 0 198 221 202
rect 585 198 630 202
rect 0 190 151 194
rect 515 190 622 194
rect 0 182 101 186
rect 465 183 614 187
rect 34 113 73 117
rect 250 114 346 117
rect 350 114 426 117
rect 370 41 373 50
rect 0 23 5 26
rect 0 18 13 23
rect 250 18 373 23
rect 605 18 640 23
rect 0 10 66 15
rect 250 10 305 15
rect 311 10 426 15
rect 610 10 640 15
rect 0 6 8 10
<< metal2 >>
rect 102 716 107 720
rect 150 719 154 720
rect 104 715 107 716
rect 148 716 154 719
rect 222 719 226 720
rect 270 719 274 720
rect 222 716 228 719
rect 148 715 152 716
rect 224 715 228 716
rect 268 716 274 719
rect 342 719 346 720
rect 390 719 394 720
rect 342 716 348 719
rect 268 715 272 716
rect 344 715 348 716
rect 388 716 394 719
rect 462 719 466 720
rect 510 719 514 720
rect 462 716 468 719
rect 388 715 392 716
rect 464 715 468 716
rect 508 716 514 719
rect 582 719 586 720
rect 582 716 588 719
rect 508 715 512 716
rect 584 715 588 716
rect 30 528 34 596
rect 30 344 34 524
rect 13 178 18 286
rect 30 117 34 340
rect 30 8 34 113
rect 38 591 42 596
rect 75 595 113 598
rect 105 593 113 595
rect 143 594 181 597
rect 195 594 233 597
rect 143 593 151 594
rect 225 591 233 594
rect 263 594 301 597
rect 315 594 353 597
rect 263 592 272 594
rect 345 591 353 594
rect 383 594 421 597
rect 435 594 473 597
rect 383 591 391 594
rect 465 592 473 594
rect 503 594 541 597
rect 555 596 572 597
rect 555 594 593 596
rect 503 592 511 594
rect 569 593 593 594
rect 569 592 581 593
rect 38 587 50 591
rect 585 590 593 593
rect 38 173 42 587
rect 75 427 79 439
rect 195 431 199 437
rect 425 430 431 437
rect 46 180 50 278
rect 66 182 71 276
rect 75 187 79 270
rect 101 266 105 270
rect 85 187 89 262
rect 125 182 131 275
rect 151 258 155 271
rect 151 186 155 190
rect 185 182 191 275
rect 195 186 199 271
rect 221 250 225 272
rect 221 186 225 198
rect 245 182 251 275
rect 271 242 275 271
rect 38 169 46 173
rect 38 0 42 169
rect 46 0 50 73
rect 305 54 311 275
rect 341 234 345 272
rect 365 184 371 276
rect 391 226 395 271
rect 365 178 378 184
rect 425 182 430 275
rect 461 218 465 271
rect 449 183 461 187
rect 485 182 491 275
rect 511 210 515 271
rect 511 183 515 190
rect 545 182 550 275
rect 581 186 585 198
rect 605 182 610 436
rect 614 187 618 643
rect 622 194 626 679
rect 630 202 634 686
rect 346 55 350 113
rect 305 50 306 54
rect 310 50 311 54
rect 305 30 311 50
rect 75 5 79 28
rect 85 11 89 29
rect 305 26 306 30
rect 310 26 311 30
rect 85 9 90 11
rect 75 2 82 5
rect 78 0 82 2
rect 86 0 90 9
rect 195 10 199 26
rect 305 15 311 26
rect 344 10 348 34
rect 195 6 202 10
rect 198 0 202 6
rect 342 7 348 10
rect 445 9 449 31
rect 342 0 346 7
rect 445 6 450 9
rect 446 0 450 6
<< m2contact >>
rect 630 686 634 690
rect 622 679 626 683
rect 614 643 618 647
rect 30 524 34 528
rect 46 479 50 483
rect 46 385 50 389
rect 30 340 34 344
rect 85 262 89 266
rect 101 262 105 266
rect 151 254 155 258
rect 221 246 225 250
rect 271 238 275 242
rect 341 230 345 234
rect 391 222 395 226
rect 461 214 465 218
rect 511 206 515 210
rect 221 198 225 202
rect 581 198 585 202
rect 630 198 634 202
rect 151 190 155 194
rect 511 190 515 194
rect 622 190 626 194
rect 101 182 105 186
rect 461 183 465 187
rect 614 183 618 187
rect 30 113 34 117
rect 346 113 350 117
rect 306 50 310 54
rect 306 26 310 30
rect 305 10 311 15
use wrapshifter wrapshifter_0
timestamp 951985653
transform 1 0 66 0 1 625
box 0 -36 544 90
use wordCounter wordCounter_0
timestamp 951112323
transform 0 -1 550 -1 0 599
box 1 -60 166 537
use pixelCounter pixelCounter_0
timestamp 951112323
transform 0 -1 130 1 0 270
box 0 -420 164 117
use pointerCounter pointerCounter_0
timestamp 951112323
transform 0 -1 253 -1 0 198
box 11 3 188 240
use countIObuffer countIObuffer_0
timestamp 951544315
transform -1 0 364 0 1 23
box -6 3 58 32
use kernelMuxCounter kernelMuxCounter_0
timestamp 951112323
transform 0 -1 505 -1 0 190
box 3 -105 180 132
<< labels >>
rlabel metal1 636 262 640 266 0 Pix_Mux_s1[7]
rlabel metal1 636 254 640 258 0 Pix_Mux_s1[6]
rlabel metal1 636 246 640 250 0 Pix_Mux_s1[5]
rlabel metal1 636 238 640 242 0 Pix_Mux_s1[4]
rlabel metal1 636 230 640 234 0 Pix_Mux_s1[3]
rlabel metal1 636 222 640 226 0 Pix_Mux_s1[2]
rlabel metal1 636 214 640 218 0 Pix_Mux_s1[1]
rlabel metal1 636 206 640 210 0 Pix_Mux_s1[0]
rlabel metal2 446 0 450 4 1 kernelCounterOut2_s1
rlabel metal1 0 6 4 10 3 Vdd
rlabel metal1 0 22 4 26 3 Gnd
rlabel metal2 38 0 42 4 1 Phi2
rlabel metal2 46 0 50 4 1 p3_Phi1_q1
rlabel metal2 78 0 82 4 1 wordCounterOut0_s1
rlabel metal2 86 0 90 4 1 pixCounterOut7_s1
rlabel metal2 198 0 202 4 1 wordCounterOut2_s1
rlabel metal2 342 0 346 4 1 Reset_s1
rlabel metal1 0 182 4 186 3 Mem_Pointer_s1[2]
rlabel metal1 0 190 4 194 3 Mem_Pointer_s1[1]
rlabel metal1 0 198 4 202 3 Mem_Pointer_s1[0]
rlabel metal1 0 478 4 482 0 c9_Phi1_q1
rlabel metal1 0 382 4 386 0 c8_Phi1_q1
rlabel metal2 102 716 106 720 0 wordCounterShifted_s1[0]
rlabel metal2 150 716 154 720 0 wordCounterShifted_s1[1]
rlabel metal2 222 716 226 720 0 wordCounterShifted_s1[2]
rlabel metal2 270 716 274 720 0 wordCounterShifted_s1[3]
rlabel metal2 342 716 346 720 0 wordCounterShifted_s1[4]
rlabel metal2 390 716 394 720 0 wordCounterShifted_s1[5]
rlabel metal2 462 716 466 720 0 wordCounterShifted_s1[6]
rlabel metal2 510 716 514 720 0 wordCounterShifted_s1[7]
rlabel metal2 582 716 586 720 0 wordCounterShifted_s1[8]
<< end >>
